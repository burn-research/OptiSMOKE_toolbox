THERMO

   300.000  1000.000  3000.000

AR                      AR  1                    298.00   3000.00 1000.00      1 ! Burcat / Goos 2016

 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2

-7.45375000E+02 4.37967491E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3

 0.00000000E+00 0.00000000E+00-7.45375000E+02 4.37967491E+00                   4

HE                      HE1                    0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2

-7.45375000E+02 9.28723974E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3

 0.00000000E+00 0.00000000E+00-7.45375000E+02 9.28723974E-01                   4

N2                      N 2                    0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2

-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3

 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00                   4

H                       H 1                    0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2

 2.54736600E+04-4.46682850E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3

 0.00000000E+00 0.00000000E+00 2.54736600E+04-4.46682850E-01                   4

O                       O 1                    0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.54363697E+00-2.73162486E-05-4.19029520E-09 4.95481845E-12-4.79553694E-16    2

 2.92260120E+04 4.92229457E+00 3.16826710E+00-3.27931884E-03 6.64306396E-06    3

-6.12806624E-09 2.11265971E-12 2.91222592E+04 2.05193346E+00                   4

OH                      H 1  O 1               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.83853033E+00 1.10741289E-03-2.94000209E-07 4.20698729E-11-2.42289890E-15    2

 3.69780808E+03 5.84494652E+00 3.99198424E+00-2.40106655E-03 4.61664033E-06    3

-3.87916306E-09 1.36319502E-12 3.36889836E+03-1.03998477E-01                   4

H2                      H 2                    0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.93286575E+00 8.26608026E-04-1.46402364E-07 1.54100414E-11-6.88804800E-16    2

-8.13065581E+02-1.02432865E+00 2.34433112E+00 7.98052075E-03-1.94781510E-05    3

 2.01572094E-08-7.37611761E-12-9.17935173E+02 6.83010238E-01                   4

O2                      O 2                    0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.66096065E+00 6.56365811E-04-1.41149627E-07 2.05797935E-11-1.29913436E-15    2

-1.21597718E+03 3.41536279E+00 3.78245636E+00-2.99673416E-03 9.84730201E-06    3

-9.68129509E-09 3.24372837E-12-1.06394356E+03 3.65767573E+00                   4

HO2                     H 1  O 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.17228741E+00 1.88117627E-03-3.46277286E-07 1.94657549E-11 1.76256905E-16    2

 3.10206839E+01 2.95767672E+00 4.30179807E+00-4.74912097E-03 2.11582905E-05    3

-2.42763914E-08 9.29225225E-12 2.64018485E+02 3.71666220E+00                   4

H2O2                    H 2  O 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.57977305E+00 4.05326003E-03-1.29844730E-06 1.98211400E-10-1.13968792E-14    2

-1.80071775E+04 6.64970694E-01 4.31515149E+00-8.47390622E-04 1.76404323E-05    3

-2.26762944E-08 9.08950158E-12-1.77067437E+04 3.27373319E+00                   4

CO                      C 1  O 1               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.04848590E+00 1.35172810E-03-4.85794050E-07 7.88536440E-11-4.69807460E-15    2

-1.42661170E+04 6.01709770E+00 3.57953350E+00-6.10353690E-04 1.01681430E-06    3

 9.07005860E-10-9.04424490E-13-1.43440860E+04 3.50840930E+00                   4

CO2                     C 1  O 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.63651110E+00 2.74145690E-03-9.95897590E-07 1.60386660E-10-9.16198570E-15    2

-4.90249040E+04-1.93489550E+00 2.35681300E+00 8.98412990E-03-7.12206320E-06    3

 2.45730080E-09-1.42885480E-13-4.83719710E+04 9.90090350E+00                   4

HCO                     C 1  H 1  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.92001542E+00 2.52279324E-03-6.71004164E-07 1.05615948E-10-7.43798261E-15    2

 3.65342928E+03 3.58077056E+00 4.23754610E+00-3.32075257E-03 1.40030264E-05    3

-1.34239995E-08 4.37416208E-12 3.87241185E+03 3.30834869E+00                   4

OH*                     H 1  O 1               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.75582920E+00 1.39848756E-03-4.19428493E-07 6.33453282E-11-3.56042218E-15    2

 5.09751756E+04 5.62581429E+00 3.46084428E+00 5.01872172E-04-2.00254474E-06    3

 3.18901984E-09-1.35451838E-12 5.07349466E+04 1.73976415E+00                   4

H2O                     H 2  O 1               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.67703890E+00 2.97318160E-03-7.73768890E-07 9.44335140E-11-4.26899910E-15    2

-2.98858940E+04 6.88255000E+00 4.19863520E+00-2.03640170E-03 6.52034160E-06    3

-5.48792690E-09 1.77196800E-12-3.02937260E+04-8.49009010E-01                   4 ! Burcat / Goos 2016

CH2O                    C 1  H 2  O 1          0300.00   3000.00  1000.00      1

 3.16952665E+00 6.19320560E-03-2.25056366E-06 3.65975660E-10-2.20149458E-14    2

-1.45486831E+04 6.04207898E+00 4.79372312E+00-9.90833322E-03 3.73219990E-05    3

-3.79285237E-08 1.31772641E-11-1.43791953E+04 6.02798058E-01                   4

CH                      C 1  H 1               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.52093690E+00 1.76536390E-03-4.61476600E-07 5.92896750E-11-3.34745010E-15    2

 7.09467690E+04 7.40518290E+00 3.48975830E+00 3.24321600E-04-1.68997510E-06    3

 3.16284200E-09-1.40618030E-12 7.06126460E+04 2.08428410E+00                   4

C                       C 1                    0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.61355965E+00-2.09502599E-04 1.13560743E-07-1.77761841E-11 9.11562299E-16    2

 8.54326029E+04 4.14774484E+00 2.55429132E+00-3.19806406E-04 7.22951974E-07    3

-7.14799930E-10 2.58116218E-13 8.54667077E+04 4.53080427E+00                   4

CH2-3                   C 1  H 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.14631886E+00 3.03671259E-03-9.96474439E-07 1.50483580E-10-8.57335515E-15    2

 4.60412605E+04 4.72341711E+00 3.71757846E+00 1.27391260E-03 2.17347251E-06    3

-3.48858500E-09 1.65208866E-12 4.58723866E+04 1.75297945E+00                   4

CH2-1                   C 1  H 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.13501686E+00 2.89593926E-03-8.16668090E-07 1.13572697E-10-6.36262835E-15    2

 5.05040504E+04 4.06030621E+00 4.19331325E+00-2.33105184E-03 8.15676451E-06    3

-6.62985981E-09 1.93233199E-12 5.03662246E+04-7.46734310E-01                   4

C2H2                    C 2  H 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.65878489E+00 4.88396667E-03-1.60828888E-06 2.46974544E-10-1.38605959E-14    2

 2.57594042E+04-3.99838194E+00 8.08679682E-01 2.33615762E-02-3.55172234E-05    3

 2.80152958E-08-8.50075165E-12 2.64289808E+04 1.39396761E+01                   4

CH3                     C 1  H 3               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 2.97812060E+00 5.79785200E-03-1.97558000E-06 3.07297900E-10-1.79174160E-14    2

 1.65095130E+04 4.72247990E+00 3.65717970E+00 2.12659790E-03 5.45838830E-06    3

-6.61810030E-09 2.46570740E-12 1.64227160E+04 1.67353540E+00                   4

CH4                     C 1  H 4               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 1.65326226E+00 1.00263099E-02-3.31661238E-06 5.36483138E-10-3.14696758E-14    2

-1.00095936E+04 9.90506283E+00 5.14911468E+00-1.36622009E-02 4.91453921E-05    3

-4.84246767E-08 1.66603441E-11-1.02465983E+04-4.63848842E+00                   4

HOCHO                   C 1  H 2  O 2          0300.00   3000.00  1000.00      1 ! Burcat / Goos 2017

 4.61383160E+00 6.44963640E-03-2.29082510E-06 3.67160470E-10-2.18736750E-14    2

-4.53303180E+04 8.47883830E-01 3.89836160E+00-3.55877950E-03 3.55205380E-05    3

-4.38499590E-08 1.71077690E-11-4.67785744E+04 7.34953970E+00                   4

CH2OH                   C 1  H 3  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.09314370E+00 5.94761260E-03-2.06497460E-06 3.23008173E-10-1.88125902E-14    2

-4.03409640E+03-1.84691493E+00 4.47834367E+00-1.35070310E-03 2.78484980E-05    3

-3.64869060E-08 1.47907450E-11-3.50072890E+03 3.30913500E+00                   4

OCHO                    C 1  H 1  O 2          0300.00   5000.00  1690.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 6.12628782E+00 3.75602932E-03-1.42010352E-06 2.36429200E-10-1.44167651E-14    2

-2.17698466E+04-8.01574694E+00 1.35213452E+00 1.50082004E-02-1.09896141E-05    3

 3.73679840E-09-4.81014498E-13-2.02253647E+04 1.74373147E+01                   4

CH3O                    C 1  H 3  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.75779238E+00 7.44142474E-03-2.69705176E-06 4.38090504E-10-2.63537098E-14    2

 3.78111940E+02-1.96680028E+00 3.71180502E+00-2.80463306E-03 3.76550971E-05    3

-4.73072089E-08 1.86588420E-11 1.29569760E+03 6.57240864E+00                   4

C2H4                    C 2  H 4               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.99182724E+00 1.04833908E-02-3.71721342E-06 5.94628366E-10-3.53630386E-14    2

 4.26865851E+03-2.69081762E-01 3.95920063E+00-7.57051373E-03 5.70989993E-05    3

-6.91588352E-08 2.69884190E-11 5.08977598E+03 4.09730213E+00                   4

CH2CO                   C 2  H 2  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.75871449E+00 6.35124053E-03-2.25955361E-06 3.62321512E-10-2.15855515E-14    2

-8.08533464E+03-4.96490444E+00 2.13241136E+00 1.81319455E-02-1.74093315E-05    3

 9.35336040E-09-2.01724844E-12-7.14808520E+03 1.33807969E+01                   4

C2H6                    C 2  H 6               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.04666411E+00 1.53538802E-02-5.47039485E-06 8.77826544E-10-5.23167531E-14    2

-1.24473499E+04-9.68698313E-01 4.29142572E+00-5.50154901E-03 5.99438458E-05    3

-7.08466469E-08 2.68685836E-11-1.15222056E+04 2.66678994E+00                   4

CH3OH                   C 1  H 4  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.52726795E+00 1.03178783E-02-3.62892944E-06 5.77448016E-10-3.42182632E-14    2

-2.60028834E+04 5.16758693E+00 5.65851051E+00-1.62983419E-02 6.91938156E-05    3

-7.58372926E-08 2.80427550E-11-2.56119736E+04-8.97330508E-01                   4

CH3O2                   C 1  H 3  O 2          0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.55530486E+00 9.12236137E-03-3.23851661E-06 5.18713798E-10-3.08834151E-14    2

-1.03569402E+03-3.99158547E+00 4.97169544E+00-5.29356557E-03 4.77334149E-05    3

-5.77065617E-08 2.22219969E-11-1.29022161E+02 2.81501182E+00                   4

CH3O2H                  C 1  H 4  O 2          0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 7.76538058E+00 8.61499712E-03-2.98006935E-06 4.68638071E-10-2.75339255E-14    2

-1.82979984E+04-1.43992663E+01 2.90540897E+00 1.74994735E-02 5.28243630E-06    3

-2.52827275E-08 1.34368212E-11-1.68894632E+04 1.13741987E+01                   4

C2H3                    C 2  H 3               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.15026763E+00 7.54021341E-03-2.62997847E-06 4.15974048E-10-2.45407509E-14    2

 3.38566380E+04 1.72812235E+00 3.36377642E+00 2.65765722E-04 2.79620704E-05    3

-3.72986942E-08 1.51590176E-11 3.44749589E+04 7.91510092E+00                   4

C2H5                    C 2  H 5               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.32195633E+00 1.23930542E-02-4.39680960E-06 7.03519917E-10-4.18435239E-14    2

 1.21759475E+04 1.71103809E-01 4.24185905E+00-3.56905235E-03 4.82667202E-05    3

-5.85401009E-08 2.25804514E-11 1.29690344E+04 4.44703782E+00                   4

C2H5OH                  C 2  H 6  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 6.56243650E+00 1.52042220E-02-5.38967950E-06 8.62250110E-10-5.12897870E-14    2

-3.15256210E+04-9.47302020E+00 4.85869570E+00-3.74017260E-03 6.95553780E-05    3

-8.86547960E-08 3.51688350E-11-2.99961320E+04 4.80185450E+00                   4

C2H5O                   C 2  H 5  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 6.55053877E+00 1.32525511E-02-4.74726060E-06 7.64699226E-10-4.57008357E-14    2

-4.47191998E+03-9.61231141E+00 3.26905655E+00 9.33562904E-03 2.96317166E-05    3

-4.53411341E-08 1.88795595E-11-2.95022955E+03 1.04200942E+01                   4

CH3CHO                  C 2  H 4  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.40411080E+00 1.17230590E-02-4.22631370E-06 6.83724510E-10-4.09848630E-14    2

-2.25931220E+04-3.48079170E+00 4.72945950E+00-3.19328580E-03 4.75349210E-05    3

-5.74586110E-08 2.19311120E-11-2.15728780E+04 4.10301590E+00                   4

CH3CO                   C 2  H 3  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.31371650E+00 9.17377930E-03-3.32203860E-06 5.39474560E-10-3.24523680E-14    2

-3.64504140E+03-1.67575580E+00 4.03587050E+00 8.77294870E-04 3.07100100E-05    3

-3.92475650E-08 1.52968690E-11-2.68207380E+03 7.86176820E+00                   4

CH2O2H                  C 1  H 3  O 2          0300.00   2500.00  1000.00      1 ! RASMUSSEN et al.; Int J Chem Kinet 40: 778â€“807, 2008

 6.98746029E+00 9.00484259E-03-3.24366912E-06 5.24324826E-10-3.13587080E-14    2

 5.01257769E+03-1.02619220E+01 5.83126679E+00-3.51771199E-03 4.54550577E-05    3

-5.66903320E-08 2.21633070E-11 6.06187060E+03-5.79143222E-01                   4

C2H                     C 2  H 1               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.66270248E+00 3.82492252E-03-1.36632500E-06 2.13455040E-10-1.23216848E-14    2

 6.71683790E+04 3.92205792E+00 2.89867676E+00 1.32988489E-02-2.80733327E-05    3

 2.89484755E-08-1.07502351E-11 6.70616050E+04 6.18547632E+00                   4

C2                      C 2                    0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 3.43350371E+00 1.07185010E-03-3.97897382E-07 6.67457391E-11-4.10152154E-15    2

 1.00178987E+05 4.10588356E+00 3.76163273E+00-2.72143299E-03 8.69879462E-06    3

-8.19304667E-09 2.62415296E-12 1.00254566E+05 3.18038623E+00                   4

C2O                     C 2  O 1               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.42468378E+00 1.85393945E-03-5.17932956E-07 6.77646230E-11-3.53315237E-15    2

 4.37161379E+04-3.69608405E+00 2.86278214E+00 1.19701204E-02-1.80851222E-05    3

 1.52777730E-08-5.20063163E-12 4.43125964E+04 8.89759099E+00                   4

HCCO                    C 2  H 1  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 5.91479333E+00 3.71408730E-03-1.30137010E-06 2.06473345E-10-1.21476759E-14    2

 1.93596301E+04-5.50567269E+00 1.87607969E+00 2.21205418E-02-3.58869325E-05    3

 3.05402541E-08-1.01281069E-11 2.01633840E+04 1.36968290E+01                   4

H2CC                    C 2  H 2               0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 4.27807305E+00 4.75622626E-03-1.63007378E-06 2.54622680E-10-1.48860086E-14    2

 4.80140478E+04 6.39978600E-01 3.28154941E+00 6.97642650E-03-2.38527914E-06    3

-1.21077631E-09 9.82041734E-13 4.83191706E+04 5.92035686E+00                   4

C3H3                    C 3  H 3               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 7.14221719E+00 7.61902211E-03-2.67460030E-06 4.24914904E-10-2.51475443E-14    2

 3.95709594E+04-1.25848690E+01 1.35110873E+00 3.27411291E-02-4.73827407E-05    3

 3.76310220E-08-1.18541128E-11 4.07679941E+04 1.52058598E+01                   4

C4H2                    C 4  H 2               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 8.68978130E+00 6.69732229E-03-2.34774865E-06 3.72759231E-10-2.20554548E-14    2

 5.19942624E+04-2.20010465E+01-5.84768273E-01 5.33506727E-02-9.50805952E-05    3

 8.37959674E-08-2.80912179E-11 5.36111160E+04 2.09878997E+01                   4

C3H5                    C 3  H 5               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2017

 6.74633155E+00 1.31071760E-02-4.60059113E-06 7.31029510E-10-4.32759674E-14    2

 1.71151431E+04-1.25248814E+01 1.65533607E+00 1.63688750E-02 2.10544223E-05    3

-4.24018394E-08 1.92638759E-11 1.89454047E+04 1.61040987E+01                   4

CH2CHO                  C 2  H 3  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 6.53928338E+00 7.80238629E-03-2.76413612E-06 4.42098906E-10-2.62954290E-14    2

-1.18858659E+03-8.72091393E+00 2.79502600E+00 1.01099472E-02 1.61750645E-05    3

-3.10303145E-08 1.39436139E-11 1.62944975E+02 1.23646657E+01                   4

C2H3OO                  C 2  H 3  O 2          0298.15   2000.00  1000.00      1 ! Aramco 2.0

 6.04483828E+00 1.45511127E-02-7.50974622E-06 1.83488280E-09-1.66689681E-13    2

 1.01699244E+04-3.71144913E+00 1.09784776E+00 2.95333237E-02-2.27744360E-05    3

 7.20559155E-09-3.07929092E-13 1.13996101E+04 2.13563583E+01                   4

HCCOH                   C 2  H 2  O 1          0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 6.37509678E+00 5.49429011E-03-1.88136576E-06 2.93803536E-10-1.71771901E-14    2

 8.93277676E+03-8.24498007E+00 2.05541154E+00 2.52003372E-02-3.80821654E-05    3

 3.09890632E-08-9.89799902E-12 9.76872113E+03 1.22271534E+01                   4

C4H4                    C 4  H 4               0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 7.98456038E+00 1.20558816E-02-4.23587475E-06 6.73646140E-10-3.99059864E-14    2

 3.11993029E+04-1.67958975E+01 1.37368786E+00 2.88801256E-02-1.46863874E-05    3

-3.91045446E-09 4.78133572E-12 3.30633344E+04 1.75941274E+01                   4

C2H2OH                  C 2  H 3  O 1          0300.00   5000.00  1401.00      1 ! Aramco 2.0

 8.20268447E+00 5.92989165E-03-1.99194448E-06 3.05794341E-10-1.76114732E-14    2

 1.24881328E+04-1.89670436E+01 6.41642616E-01 2.61903633E-02-2.30385370E-05    3

 1.02804704E-08-1.81971416E-12 1.48276951E+04 2.06750999E+01                   4

C2H3CHO                 C 3  H 4  O 1          0298.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 8.20654919E+00 1.28492916E-02-4.64285331E-06 7.51738738E-10-4.51298116E-14    2

-1.18838341E+04-1.49881933E+01 4.69868861E+00 4.99965957E-03 4.38587397E-05    3

-6.12883900E-08 2.48508985E-11-1.00875286E+04 7.29812046E+00                   4

C3H4O                   C 3  H 4  O 1          0300.00   3000.00  1000.00      1 ! Seidel et al. 2015 cited Burcat / Goos 2016

 8.20654919E+00 1.28492916E-02-4.64285331E-06 7.51738738E-10-4.51298116E-14    2

-1.18838341E+04-1.49881933E+01 4.69868861E+00 4.99965957E-03 4.38587397E-05    3

-6.12883900E-08 2.48508985E-11-1.00875286E+04 7.29812046E+00                   4

CHCHO                   C 2  H 2  O 1          0298.15   2000.00  1000.00      1 ! Aramco 2.0

 4.92632910E+00 9.71712147E-03-5.54855980E-06 1.53068537E-09-1.64742462E-13    2

 2.89499494E+04 5.27874677E-01 2.33256751E+00 1.62952986E-02-9.72052177E-06    3

 5.15124155E-10 1.03836514E-12 2.96585452E+04 1.39904923E+01                   4

CHOCHO                  C 2  H 2  O 2          0300.00   5000.00  1386.00      1 ! Aramco 2.0

 9.75438561E+00 4.97645947E-03-1.74410483E-06 2.75586994E-10-1.61969892E-14    2

-2.95832896E+04-2.61878329E+01 1.88105120E+00 2.36386368E-02-1.83443295E-05    3

 6.84842963E-09-9.92733674E-13-2.69280190E+04 1.59154793E+01                   4

CHOCO                   C 2  H 1  O 2          0300.00   5000.00  1000.00      1 ! Togbe et al. 2011; PROCI 33 (2011) 367â€“374

 8.35919700E+00 4.49470900E-03-1.98795700E-06 3.89038900E-10-2.79353800E-14    2

-1.24067300E+04-1.67672000E+01 7.66973900E+00-1.29080300E-02 5.95280900E-05    3

-6.96004300E-08 2.65376800E-11-1.13370100E+04-8.67146000E+00                   4

CH3CO2                  C 2  H 3  O 2          0300.00   3000.00  1000.00      1 ! Burcat / Goos 2016

 7.62274600E+00 9.66664529E-03-3.47122481E-06 5.60301057E-10-3.35405698E-14    2

-2.63946612E+04-1.31344143E+01 2.81652185E+00 1.74597055E-02 1.83449161E-06    3

-1.54957310E-08 7.72993893E-12-2.47922272E+04 1.30310283E+01                   4

CH3CO3                  C 2  H 3  O 3          0300.00   3000.00  1391.00      1 ! Seidel et al. 2015;

 1.12522498E+01 8.33652672E-03-2.89014530E-06 4.52781734E-10-2.64354456E-14    2

-2.60238584E+04-2.96370457E+01 3.60373432E+00 2.70080341E-02-2.08293438E-05    3

 8.50541104E-09-1.43846110E-12-2.34205171E+04 1.12014914E+01                   4

CH3CO3H                 C 2  H 4  O 3          0300.00   3000.00  1391.00      1 ! Seidel et al. 2015;

 1.25060485E+01 9.47789695E-03-3.30402246E-06 5.19630793E-10-3.04233568E-14    2

-4.59856703E+04-3.79195947E+01 2.24135876E+00 3.37963514E-02-2.53887482E-05    3

 9.67583587E-09-1.49266157E-12-4.24677831E+04 1.70668133E+01                   4

C3H6                    C 3  H 6               0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 6.03870234E+00 1.62963931E-02-5.82130800E-06 9.35936829E-10-5.58603143E-14    2

-7.41715057E+02-8.43825992E+00 3.83464468E+00 3.29078952E-03 5.05228001E-05    3

-6.66251176E-08 2.63707473E-11 7.88717123E+02 7.53408013E+00                   4

C3H8                    C 3  H 8               0298.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 6.66919760E+00 2.06108751E-02-7.36512349E-06 1.18434262E-09-7.06914630E-14    2

-1.62754066E+04-1.31943379E+01 4.21093013E+00 1.70886504E-03 7.06530164E-05    3

-9.20060565E-08 3.64618453E-11-1.43810883E+04 5.61004451E+00                   4

I-C3H7                  C 3  H 7               0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 5.30597255E+00 1.89854588E-02-6.74315384E-06 1.07993730E-09-6.42785036E-14    2

 7.78748910E+03-2.23233935E+00 5.47421257E+00-8.42536682E-03 8.04607759E-05    3

-9.49287824E-08 3.59830971E-11 9.04939013E+03 3.40542323E+00                   4

N-C3H7                  C 3  H 7               0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 6.49636579E+00 1.77337992E-02-6.24898046E-06 9.95389495E-10-5.90199770E-14    2

 8.85973885E+03-8.56389710E+00 4.08211458E+00 5.23240341E-03 5.13554466E-05    3

-6.99343598E-08 2.81819493E-11 1.04074558E+04 8.39534919E+00                   4

C3H4                    C 3  H 4               0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 6.31687220E+00 1.11337280E-02-3.96293780E-06 6.35642380E-10-3.78755400E-14    2

 2.01174950E+04-1.09957660E+01 2.61304450E+00 1.21225750E-02 1.85398800E-05    3

-3.45251490E-08 1.53350790E-11 2.15415670E+04 1.02261390E+01                   4

C3H4P                   C 3  H 4               0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 6.02524000E+00 1.13365420E-02-4.02233910E-06 6.43760630E-10-3.82996350E-14    2

 1.96209420E+04-8.60437850E+00 2.68038690E+00 1.57996510E-02 2.50705960E-06    3

-1.36576230E-08 6.61542850E-12 2.08023740E+04 9.87693510E+00                   4

CH2CHOH                 C 2  H 4  O 1          0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 7.20200781E+00 9.59749604E-03-3.34348031E-06 5.28604398E-10-3.11832760E-14    2

-1.79990363E+04-1.34267646E+01 1.95966153E+00 2.01744811E-02-1.09658218E-06    3

-1.62414813E-08 9.15736550E-12-1.64393370E+04 1.43785378E+01                   4

CH3CHOH                 C 2  H 5  O 1          0298.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 6.35842302E+00 1.24356276E-02-4.33096839E-06 6.84530381E-10-4.03713238E-14    2

-9.53018581E+03-6.05106112E+00 4.22283250E+00 5.12174798E-03 3.48386522E-05    3

-4.91943637E-08 2.01183723E-11-8.35622088E+03 8.01675700E+00                   4

CH2CH2OH                C 2  H 5  O 1          0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2017 

 7.01348674E+00 1.20204391E-02-4.21992012E-06 6.70675981E-10-3.97135273E-14    2

-6.16161779E+03-8.62052409E+00 4.20954137E+00 9.12964578E-03 2.47462263E-05    3

-3.92945764E-08 1.66541312E-11-4.91511371E+03 8.30445413E+00                   4

C2H5O2                  C 2  H 5  O 2          0300.00   5000.00  1389.00      1 ! Burke et al. 2014;  Combustion and Flame 161 (2014) 2765â€“2784

 9.50282570E+00 1.20429839E-02-4.09491581E-06 6.33049241E-10-3.66133788E-14    2

-7.37069391E+03-2.21717130E+01 3.90351912E+00 2.22599212E-02-1.01610079E-05    3

 1.71709751E-09 1.88166738E-14-5.09654081E+03 8.98722750E+00                   4

C2H4O1-2                C 2  H 4  O 1          0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 5.48876410E+00 1.20461900E-02-4.33369310E-06 7.00283110E-10-4.19490880E-14    2

-9.18042510E+03-7.07996050E+00 3.75905320E+00-9.44121800E-03 8.03097210E-05    3

-1.00807880E-07 4.00399210E-11-7.56081430E+03 7.84974750E+00                   4

C2H5O2H                 C 2  H 6  O 2          0298.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 9.58691079E+00 1.48603589E-02-5.29787964E-06 8.47317148E-10-5.03436325E-14    2

-2.38367900E+04-2.28310676E+01 4.14672004E+00 9.78668137E-03 4.91492257E-05    3

-7.42532076E-08 3.11169441E-11-2.14671219E+04 9.84024999E+00                   4

C2H5CHO                 C 3  H 6  O 1          0298.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 7.44085690E+00 1.77301764E-02-6.34081568E-06 1.02040803E-09-6.09461714E-14    2

-2.60055814E+04-1.44195446E+01 4.24529681E+00 6.68296706E-03 4.93337933E-05    3

-6.71986124E-08 2.67262347E-11-2.41473007E+04 6.90738560E+00                   4

C2H5CO                  C 3  H 5  O 1          0298.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 6.52325448E+00 1.54211952E-02-5.50898157E-06 8.85889862E-10-5.28846399E-14    2

-7.19631634E+03-5.19862218E+00 6.25722402E+00-9.17612184E-03 7.61190493E-05    3

-9.05514997E-08 3.46198215E-11-5.91616484E+03 2.23330599E+00                   4

C2H4O2H                 C 2  H 5  O 2          0300.00   5000.00  1389.00      1 ! Burke et al. 2014;  Combustion and Flame 161 (2014) 2765â€“2784

 1.00590614E+01 1.13378955E-02-3.89403387E-06 6.06090687E-10-3.52212353E-14    2

 4.24048653E+02-2.32086536E+01 2.75788364E+00 2.88271987E-02-2.08302264E-05    3

 8.47401397E-09-1.48617610E-12 3.00153893E+03 1.59921711E+01                   4

C2H3O1-2                C 2  H 3  O 1          0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 5.60158035E+00 9.17613962E-03-3.28028902E-06 5.27903888E-10-3.15362241E-14    2

 1.71446252E+04-5.47228512E+00 3.58349017E+00-6.02275805E-03 6.32426867E-05    3

-8.18540707E-08 3.30444505E-11 1.85681353E+04 9.59725926E+00                   4

CH3OCH3-DME             C 2  H 6  O 1          0300.00   3000.00  1000.00      1 ! Burcat/ Goos 2016

 5.64844274E+00 1.63381875E-02-5.86802189E-06 9.46836384E-10-5.66504295E-14    2

-2.50864216E+04-5.96267354E+00 5.30562273E+00-2.14253958E-03 5.30873092E-05    3

-6.23146897E-08 2.30730916E-11-2.39655820E+04 7.13244569E-01                   4

CH3OCH2                 C 2  H 5  O 1          0300.00   5000.00  1376.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 8.17137842E+00 1.10086181E-02-3.82352277E-06 5.99637202E-10-3.50317513E-14    2

-3.41941605E+03-1.78650856E+01 2.91327415E+00 2.03364659E-02-9.59712342E-06    3

 2.07478525E-09-1.71343362E-13-1.18844240E+03 1.16066817E+01                   4

CH3OCH2O2               C 2  H 5  O 3          0300.00   5000.00  1389.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.24249729E+01 1.18705986E-02-4.07906532E-06 6.35310809E-10-3.69427867E-14    2

-2.29679238E+04-3.53740145E+01 2.21029612E+00 3.68877454E-02-2.82561555E-05    3

 1.15730533E-08-1.97130470E-12-1.94940940E+04 1.91463601E+01                   4

CH3OCH2O2H              C 2  H 6  O 3          0300.00   5000.00  1392.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.49370964E+01 1.19465829E-02-4.12746359E-06 6.45422590E-10-3.76427939E-14    2

-4.11001068E+04-4.99552737E+01 1.19855761E+00 4.59060764E-02-3.66252420E-05    3

 1.49318970E-08-2.46057445E-12-3.65363161E+04 2.31339904E+01                   4

CH3OCH2O                C 2  H 5  O 2          0300.00   5000.00  2012.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 8.60261845E+00 1.35772195E-02-4.84661602E-06 7.77766193E-10-4.62633624E-14    2

-2.13762444E+04-1.75775023E+01 3.25889339E+00 2.22146359E-02-7.78556340E-06    3

-2.41484158E-10 4.51914496E-13-1.92377212E+04 1.23680069E+01                   4

CH3OCHO                 C 2  H 4  O 2          0300.00   5000.00  1686.00      1 ! Zhao 2008;; Int J Chem Kinet 40: 1â€“18, 2008 

 8.69123518E+00 1.15503122E-02-4.27782486E-06 7.02533059E-10-4.24333552E-14    2

-4.64364769E+04-1.89301478E+01 3.08839783E+00 2.03760048E-02-6.84777040E-06    3

-7.28186203E-10 5.62130216E-13-4.41855167E+04 1.25364719E+01                   4

CH2OCHO                 C 2  H 3  O 2          0300.00   5000.00  1442.00      1 ! Burke 2015;Combustion and Flame 162 (2015) 315â€“330

 1.00960096E+01 7.19887066E-03-2.59813465E-06 4.18110812E-10-2.48723387E-14    2

-2.36389018E+04-2.71144175E+01 2.31031671E+00 1.80474065E-02-2.71519637E-06    3

-4.60918579E-09 1.70037078E-12-2.02910878E+04 1.71549722E+01                   4

CH3OCO                  C 2  H 3  O 2          0300.00   5000.00  1362.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.30877600E+01 4.53544950E-03-1.65096364E-06 2.67197277E-10-1.59576863E-14    2

-2.46616400E+04-3.27914051E+01 3.94199159E+00 2.43434884E-02-1.65595560E-05    3

 4.58537411E-09-3.31795708E-13-2.14404829E+04 1.66954362E+01                   4

CH2OCH2O2H              C 2  H 5  O 3          0300.00   5000.00  1393.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.51191783E+01 9.23718883E-03-3.19127505E-06 4.99114678E-10-2.91162488E-14    2

-1.84114867E+04-4.85706618E+01 2.52895507E+00 4.24128290E-02-3.73406386E-05    3

 1.66639333E-08-2.96443312E-12-1.44293306E+04 1.76899251E+01                   4

O2CH2OCH2O2H            C 2  H 5  O 5          0300.00   5000.00  1402.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.92038046E+01 1.04394841E-02-3.60582939E-06 5.63792843E-10-3.28807214E-14    2

-3.79207055E+04-6.51847273E+01 1.99640551E+00 5.83226232E-02-5.53259778E-05    3

 2.59810540E-08-4.77141005E-12-3.27628742E+04 2.44215005E+01                   4

HO2CH2OCHO              C 2  H 4  O 4          0300.00   5000.00  1387.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.64584298E+01 8.52683511E-03-3.04113500E-06 4.85596908E-10-2.87316334E-14    2

-6.23959608E+04-5.38924139E+01 3.47935703E+00 4.02952392E-02-3.30109296E-05    3

 1.34360117E-08-2.18601580E-12-5.80629934E+04 1.52521392E+01                   4

OCH2OCHO                C 2  H 3  O 3          0300.00   5000.00  1475.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.20233916E+01 8.11262659E-03-2.91356462E-06 4.67340384E-10-2.77375525E-14    2

-4.33647231E+04-3.33691809E+01 5.19690837E+00 1.58839723E-02 3.53540547E-07    3

-6.10456923E-09 1.94661801E-12-4.02242792E+04 6.11645828E+00                   4

HOCH2OCO                C 2  H 3  O 3          0300.00   5000.00  1603.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 1.13737391E+01 8.17663898E-03-2.92034021E-06 4.66695616E-10-2.76276823E-14    2

-4.65575743E+04-2.86035265E+01 6.08180801E+00 1.28768359E-02 2.04419418E-06    3

-6.10154921E-09 1.79820559E-12-4.39526183E+04 2.54054449E+00                   4

HOCH2O                  C 1  H 3  O 2          0300.00   5000.00  1452.00      1 ! Zhao 2008; Int J Chem Kinet 40: 1â€“18, 2008

 6.39521515E+00 7.43673043E-03-2.50422354E-06 3.84879712E-10-2.21778689E-14    2

-2.47500385E+04-7.29290847E+00 4.11183145E+00 7.53850697E-03 3.77337370E-06    3

-5.38746005E-09 1.45615887E-12-2.34414546E+04 6.81381989E+00                   4

CH*                     C 1  H 1               0298.00   3000.00  1000.00      1 ! Burcat/Goos 2016

 2.78220752E+00 1.47246754E-03-4.63436227E-07 7.32736021E-11-4.19705404E-15    2

 1.04547060E+05 5.17421018E+00 3.47250101E+00 4.26443626E-04-1.95181794E-06    3

 3.51755043E-09-1.60436174E-12 1.04334869E+05 1.44799533E+00                   4

!---------------NOx Thermo data starts here------------------------------------

!Thermodata for NOx Chemistry from Lamoureux 2016 taken from this very work

!for the species that are in their mechanism; additional species included in this

!mechanism are adopted from Burcat thermochemistry data base and for other sources

!see the comment

HCN               ATcT/AH  1.C  1.N  1.   0.G   200.000  6000.000 1000.00      1 ! Lamoureux et al. 2016

 3.80231648E+00 3.14630087E-03-1.06315727E-06 1.66185438E-10-9.79891962E-15    2

 1.42849502E+04 1.57501632E+00 2.25901199E+00 1.00510475E-02-1.33514567E-05    3

 1.00920479E-08-3.00880408E-12 1.45903166E+04 8.91631960E+00 1.56111424E+04    4

HCNO Fulminic AcidA 5/05H  1.N  1.C  1.O  1.G   200.000  6000.000 1000.00      1 ! Lamoureux et al. 2016

 5.91979744E+00 4.00114600E-03-1.42063343E-06 2.27569621E-10-1.35504870E-14    2

 1.80385534E+04-8.26935223E+00 6.07949401E-01 2.82182431E-02-4.60451618E-05    3

 3.82559486E-08-1.23226501E-11 1.90714209E+04 1.69199098E+01 2.01698706E+04    4

HNC               ATcT/AH  1.N  1.C  1.   0.G   200.000  6000.000 1000.00      1 ! Lamoureux et al. 2016

 4.22248262E+00 2.59458082E-03-8.58480324E-07 1.30744940E-10-7.50339813E-15    2

 2.17156730E+04-7.79706410E-02 2.30186822E+00 1.54157449E-02-3.13261898E-05    3

 3.08816218E-08-1.11912204E-11 2.19306327E+04 8.14749128E+00 2.30810956E+04    4

HNCN Cyanamide    T03/10C  1.H  1.N  2.   0.G   200.000  6000.000 1000.        1 ! Lamoureux et al. 2016

 5.53846448E+00 3.89054126E-03-1.38104752E-06 2.21294765E-10-1.31827325E-14    2

 3.59635337E+04-3.39587098E+00 3.06754311E+00 1.06789939E-02-7.96224305E-06    3

 2.59883390E-09-1.27057612E-13 3.66623508E+04 9.41074995E+00 3.79863165E+04    4

HNCO Isocyanic AciA 5/05H  1.N  1.C  1.O  1.G   200.000  6000.000 1000.00      1 ! Lamoureux et al. 2016

 5.30045051E+00 4.02250821E-03-1.40962280E-06 2.23855342E-10-1.32499966E-14    2

-1.61995274E+04-3.11770684E+00 2.24009031E+00 1.45600497E-02-1.54352330E-05    3

 8.55535028E-09-1.79631611E-12-1.54589951E+04 1.21663775E+01-1.42642740E+04    4

HNO               121286H   1N   1O   1     G  0300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.03615144E+02 0.03212486E-01-0.01260337E-04 0.02267298E-08-0.01536236E-12    2

 0.01066191E+06 0.04810264E+02 0.02784403E+02 0.06609646E-01-0.09300223E-04    3

 0.09437980E-07-0.03753146E-10 0.01091878E+06 0.09035629E+02                   4

!HNO                     H   1N   1O   1     G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 2.58819802E+00 4.87708822E-03-2.29243315E-06 5.82214028E-10-5.94811743E-14    2

! 1.20213574E+04 1.04315796E+01 4.51988078E+00-5.42507623E-03 1.70239636E-05    3

!-1.48708172E-08 4.44763498E-12 1.17637925E+04 1.75618526E+00                   4

HOCN Cyanic Acid  A 5/05H  1.N  1.C  1.O  1.G   200.000  6000.000 1000.0       1 ! Lamoureux et al. 2016

 5.28767714E+00 4.01746511E-03-1.40407465E-06 2.22562614E-10-1.31562375E-14    2

-3.77409807E+03-2.64470976E+00 2.88943546E+00 1.16487242E-02-1.08005006E-05    3

 5.44138776E-09-1.06857286E-12-3.15296691E+03 9.51295652E+00-1.85890558E+03    4

HONO               31787H   1N   1O   2     G  0300.00   5000.00  1000.00      1 ! Nitrous acid  ! Lamoureux et al. 2016

 0.05486893E+02 0.04218065E-01-0.01649143E-04 0.02971877E-08-0.02021148E-12    2 ! Also used by Dayma 2007; PROCI 31 (2007) 411â€“418

-0.01126865E+06-0.02997002E+02 0.02290413E+02 0.01409922E+00-0.01367872E-03    3

 0.07498780E-07-0.01876905E-10-0.01043195E+06 0.01328077E+03                   4

!HONO                    H   1N   1O   2     G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 4.19966671E+00 5.94217338E-03-2.95404834E-06 7.19846187E-10-6.74909061E-14    2 ! it is HONOtrans 

!-1.08122769E+04 5.08809833E+00 3.49106617E+00 6.81116875E-03-1.30943120E-06    3

!-2.34197204E-09 1.18931535E-12-1.05722865E+04 8.99803804E+00                   4

!HONO trans  Nitrous acid  SIGMA=1  STATWT=1  IA=0.9077  IB=6.681  IC=7.5887   

!Nu=3703,1795,1324,864,630.5,596  REF=Burcat G3B3  HF298=-79.190+/-0.077 kJ

!REF=Ruscic ATcT D 2013  {HF298=-79.617+/-8. kJ  REF=Burcat G3B3}  Max Lst Sq

!Error Cp @ 6000 K 0.31%.

!HONO  trans       T 2/14H  1.N  1.O  2.   0.G   200.000  6000.000  1000.00     1 ! Burcat 2017

! 5.59069580E+00 3.76633148E-03-1.32079549E-06 2.10072062E-10-1.24546207E-14    2 !

!-1.16009741E+04-3.66793086E+00 2.55834541E+00 1.11295585E-02-5.09304078E-06    3 !

!-2.76314117E-09 2.40212731E-12-1.07324351E+04 1.21891248E+01-9.52431352E+03    4 !

N                 120186N   1               G  0300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.02450268E+02 0.01066146E-02-0.07465337E-06 0.01879652E-09-0.01025984E-13    2

 0.05611604E+06 0.04448758E+02 0.02503071E+02-0.02180018E-03 0.05420529E-06    3

-0.05647560E-09 0.02099904E-12 0.05609890E+06 0.04167566E+02                   4

H2NO              102290H   2N   1O   1     G  0300.00   4000.00  1500.00      1 ! Lamoureux et al. 2016

 0.05673346E+02 0.02298837E-01-0.01774446E-05-0.01103482E-08 0.01859762E-12    2

 0.05569325E+05-0.06153540E+02 0.02530590E+02 0.08596035E-01-0.05471030E-04    3

 0.02276249E-07-0.04648073E-11 0.06868030E+05 0.01126651E+03                   4

H2CN               41687H   2C   1N   1     G  0300.00   4000.00  1000.00      1 ! Lamoureux et al. 2016

 0.05209703E+02 0.02969291E-01-0.02855589E-05-0.01635550E-08 0.03043259E-12    2

 0.02767711E+06-0.04444478E+02 0.02851661E+02 0.05695233E-01 0.01071140E-04    3

-0.01622612E-07-0.02351108E-11 0.02863782E+06 0.08992751E+02                   4

N2H2              121286N   2H   2          G  0300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.03371185E+02 0.06039968E-01-0.02303854E-04 0.04062789E-08-0.02713144E-12    2

 0.02418172E+06 0.04980585E+02 0.01617999E+02 0.01306312E+00-0.01715712E-03    3

 0.01605608E-06-0.06093639E-10 0.02467526E+06 0.01379467E+03                   4

N2O               121286N   2O   1          G   300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.04718977E+02 0.02873714E-01-0.01197496E-04 0.02250552E-08-0.01575337E-12    2

 0.08165811E+05-0.01657250E+02 0.02543058E+02 0.09492193E-01-0.09792775E-04    3

 0.06263845E-07-0.01901826E-10 0.08765100E+05 0.09511222E+02                   4

!NCN GOOS+Friedric T 1/12N   2C   1   0     0G   200.000  6000.000 1000.00      1 ! Lamoureux 2016 : adjusted a6 term which is mentioned in there paper

! 5.68743460E+00 1.82663439E-03-7.07551130E-07 1.19517763E-10-7.31862017E-15    2

! 5.14021222E+04-6.31950475E+00 2.79807986E+00 1.00008861E-02-9.59242059E-06    3

! 4.75565678E-09-1.04348512E-12 5.22141728E+04 8.62129570E+00 5.50603704E+04    4

NCN                     N   2C  1.   0.    0G   200.000  6000.000 1000.00      1 !  Goos et.al. 2013; PROCI 34 (2013) 657â€“666

 5.68743460E+00 1.82663439E-03-7.07551130E-07 1.19517763E-10-7.31862017E-15    2 !

 5.30454071E+04-6.31950475E+00 2.79807986E+00 1.00008861E-02-9.59242059E-06    3 !

 4.75565678E-09-1.04348512E-12 5.38574577E+04 8.62129570E+00 5.50603704E+04    4 !

!NCN  MethaneTetr        N   2C  1.   0.    0G   200.000  6000.000 1000.00      1 ! Burcat 2017 : REF=JACOX JPCRD (1998) & GURVICH 91

! 5.68744173E+00 1.82662756E-03-7.07546249E-07 1.19515592E-10-7.31827071E-15    2 ! HF298=445.73+/-1.7 kJ   REF=ATcT C

! 5.15901177E+04-6.31954433E+00 2.79807977E+00 1.00008683E-02-9.59229469E-06    3 ! E.Goos et al Proc Comb Symp 2012;

! 4.75546842E-09-1.04340146E-12 5.24021705E+04 8.62129767E+00 5.36050832E+04    4 ! Max Lst Sq Error Cp @ 1300 K 0.36%.

!NCN                     C   1N   2          G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 4.47903710E+00 4.18411508E-03-2.63288979E-06 7.49201653E-10-8.04623880E-14    2 ! HF298=454.57+/-1.8 kJ

! 5.30622825E+04 1.83947963E-01 3.15727170E+00 7.25557223E-03-3.91666888E-06    3 !

!-6.10550047E-10 8.13376644E-13 5.34374158E+04 7.11460304E+00                   4 !

NCO  (CNO)        A 5/05N  1.C  1.O  1.   0.G   200.000  6000.000 1000.00      1  ! Lamoureux et al. 2016

 5.08064474E+00 2.37443587E-03-9.07098904E-07 1.52286713E-10-9.31009234E-15    2

 1.35781204E+04-2.15734434E+00 2.77405177E+00 9.24523481E-03-9.91773586E-06    3

 6.68461303E-09-2.09520542E-12 1.42369570E+04 9.75458670E+00 1.53995606E+04    4

NH                 31387H   1N   1          G  0300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.02760249E+02 0.01375346E-01-0.04451914E-05 0.07692792E-09-0.05017592E-13    2

 0.04207828E+06 0.05857199E+02 0.03339758E+02 0.01253009E-01-0.03491646E-04    3

 0.04218812E-07-0.01557618E-10 0.04185047E+06 0.02507181E+02                   4

!NH                      H   1N   1          G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 2.95100955E+00 9.09994439E-04-8.35582439E-08-5.17312027E-11 1.13981436E-14    2

! 4.19707045E+04 4.83056694E+00 3.44697209E+00 5.57847818E-04-2.00289360E-06    3

! 2.85952922E-09-1.12434284E-12 4.17899268E+04 2.02990852E+00                   4

NH2               121686N   1H   2          G  0300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.02961311E+02 0.02932699E-01-0.09063600E-05 0.01617257E-08-0.01204200E-12    2

 0.02191977E+06 0.05777878E+02 0.03432493E+02 0.03299540E-01-0.06613600E-04    3

 0.08590947E-07-0.03572047E-10 0.02177228E+06 0.03090111E+02                   4

!NH2                     H   2N   1          G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 2.62839610E+00 3.44379888E-03-1.08606365E-06 1.50714038E-10-4.59423280E-15    2

! 2.15909586E+04 7.65372613E+00 3.97883538E+00-5.13888088E-04 2.68436156E-06    3

!-9.18832600E-10-9.82251152E-14 2.12486673E+04 7.77619668E-01                   4

!NH2           RAD IU3/03N   1H   2          G  0300.00   5000.00  1000.00      1 ! Burcat 2017

! 2.59263049E+00 3.47683597E-03-1.08271624E-06 1.49342558E-10-5.75241187E-15    2

! 2.18865421E+04 7.90565351E+00 4.19198016E+00-2.04602827E-03 6.67756134E-06    3

!-5.24907235E-09 1.55589948E-12 2.14991387E+04-9.04785244E-02 2.27072912E+04    4

NH3               121386N   1H   3          G  0300.00   5000.00  1000.00      1 ! Lamoureux 2016

 0.02461904E+02 0.06059166E-01-0.02004977E-04 0.03136003E-08-0.01938317E-12    2

-0.06493270E+05 0.07472097E+02 0.02204352E+02 0.01011476E+00-0.01465265E-03    3

 0.01447235E-06-0.05328509E-10-0.06525488E+05 0.08127138E+02                   4

!NH3                     H   3N   1          G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 1.07096958E+00 8.75466951E-03-3.33525419E-06 4.72015791E-10-1.13562571E-14    2

!-5.77168689E+03 1.49517392E+01 3.26650510E+00 3.05892867E-03 5.78755223E-07    3

! 9.49077412E-10-9.02221969E-13-6.36511405E+03 3.58794921E+00                   4

NNH               T 8/11N  2.H  1.   0.   0.G   200.000  6000.000 1000.00      1 ! Lamoureux et al. 2016

 3.42744423E+00 3.23295234E-03-1.17296299E-06 1.90508356E-10-1.14491506E-14    2

 2.87676026E+04 6.39209233E+00 4.25474632E+00-3.45098298E-03 1.37788699E-05    3

-1.33263744E-08 4.41023397E-12 2.87932080E+04 3.28551762E+00 3.00058572E+04    4

NO                121286N   1O   1          G   300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.03245435E+02 0.01269138E-01-0.05015890E-05 0.09169283E-09-0.06275419E-13    2

 0.09800840E+05 0.06417294E+02 0.03376542E+02 0.01253063E-01-0.03302751E-04    3

 0.05217810E-07-0.02446263E-10 0.09817961E+05 0.05829590E+02                   4

NO2               121286N   1O   2          G   300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.04682859E+02 0.02462429E-01-0.01042259E-04 0.01976902E-08-0.01391717E-12    2

 0.02261292E+05 0.09885985E+01 0.02670600E+02 0.07838501E-01-0.08063865E-04    3

 0.06161715E-07-0.02320150E-10 0.02896291E+05 0.01161207E+03                   4

!NO                      N   1O   1          G   298.150  3000.000 1000.00      1 ! Bugler 2016

! 2.79462839E+00 2.12260586E-03-1.11936971E-06 2.79521018E-10-2.68625363E-14    2

! 1.00019069E+04 8.88322674E+00 4.15036687E+00-4.08890008E-03 9.38071726E-06    3

!-7.50908901E-09 2.11742798E-12 9.77018679E+03 2.53971032E+00                   4

!NO2                     N   1O   2          G   298.150  3000.000 1000.00      1 ! Bugler 2016

! 3.65239279E+00 4.71632310E-03-2.74591748E-06 7.45382834E-10-7.63891108E-14    2

! 2.57216137E+03 6.52683440E+00 3.39100918E+00 2.62448348E-03 5.09790306E-06    3

!-7.62120493E-09 2.79960135E-12 2.78130679E+03 8.57220275E+00                   4

C2N2                    C   2N   20   00   0G   300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

 0.65480000E+01 0.39847100E-02-0.16342200E-05 0.30386000E-09-0.21110000E-13    2

 0.34907200E+05-0.97360000E+01 0.42654600E+01 0.11922570E-01-0.13420140E-04    3

 0.91923000E-08-0.27789400E-11 0.35478900E+05 0.17130000E+01                   4

HCNN              SRI/94C   1N   2H   1     G   300.000  5000.000  1000.000    1 ! Lamoureux et al. 2016

 0.58946362E+01 0.39895959E-02-0.15982380E-05 0.29249395E-09-0.20094686E-13    2

 0.53452941E+05-0.51030502E+01 0.25243194E+01 0.15960619E-01-0.18816354E-04    3

 0.12125540E-07-0.32357378E-11 0.54261984E+05 0.11675870E+02                   4

!CN   Canneaux     060110C   1N   1          G  0300.00   5000.00  1000.00      1 ! Lamoureux et al. 2016

! 3.07579471E+00 1.39061179E-03-5.54920326E-07 1.00883206E-10-6.88175427E-15    2

! 5.24171303E+04 6.38512235E+00 3.52489264E+00-2.57015392E-04 2.11721936E-07    3

! 1.77403167E-09-1.26029239E-12 5.23686935E+04 4.30280631E+00                   4

CN                IU8/03C   1N   1         0G    200.00   6000.00 1000.0       1 ! E. Goos, A. Burcat, and B. Ruscic

 3.39912850E+00 7.46548662E-04-1.41493852E-07 1.86747736E-11-1.26032540E-15    2 ! Accessed 2018

 5.16569715E+04 4.67148681E+00 3.61256069E+00-9.53015737E-04 2.13757271E-06    3

-3.05001808E-10-4.70518097E-13 5.17084034E+04 3.98238722E+00 5.27611901E+04    4

N2H3  Hydrazine   A05/05H  3.N  2.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat/Goos 2017

 4.04483566E+00 7.31130186E-03-2.47625799E-06 3.83733021E-10-2.23107573E-14    2

 2.48098603E+04 2.88423392E+00 3.42125505E+00 1.34901590E-03 2.23459071E-05    3

-2.99727732E-08 1.20978970E-11 2.53056139E+04 7.83176309E+00 2.65295249E+04    4

N2H4 HYDRAZINE    L 5/90N   2H   4    0    0G   200.000  6000.000 1000.00      1 ! Burcat/Goos 2017

 4.93957357E+00 8.75017187E-03-2.99399058E-06 4.67278418E-10-2.73068599E-14    2

 9.28265548E+03-2.69439772E+00 3.83472149E+00-6.49129555E-04 3.76848463E-05    3

-5.00709182E-08 2.03362064E-11 1.00893925E+04 5.75272030E+00 1.14474575E+04    4

H2NN Isodiazene   T 9/11N  2.H  2.   0.   0.G   200.000  6000.000  1000.00     1 ! Burcat/Goos 2017

 3.05903670E+00 6.18382347E-03-2.22171165E-06 3.58539206E-10-2.14532905E-14    2

 3.48530149E+04 6.69893515E+00 4.53204001E+00-7.32418578E-03 3.00803713E-05    3

-3.04000551E-08 1.04700639E-11 3.49580003E+04 1.51074195E+00 3.61943157E+04    4

HNOH trans & Equ  T11/11H  2.N  1.O  1.   0.G   200.000  6000.000  1000.00     1 ! Burcat/Goos 2017

 3.98321933E+00 4.88846374E-03-1.65086637E-06 2.55371446E-10-1.48308561E-14    2

 1.05780106E+04 3.62582838E+00 3.95608248E+00-3.02611020E-03 2.56874396E-05    3

-3.15645120E-08 1.24084574E-11 1.09199790E+04 5.55950983E+00 1.21354115E+04    4

NH2OH             ATcT/AN  1.H  3.O  1.   0.G   200.000  6000.000 1000.0       1 ! Burcat/Goos 2017

 3.88112502E+00 8.15708448E-03-2.82615576E-06 4.37930933E-10-2.52724604E-14    2

-6.86018419E+03 3.79156136E+00 3.21016092E+00 6.19671676E-03 1.10594948E-05    3

-1.96668262E-08 8.82516590E-12-6.58148481E+03 7.93293571E+00-5.28593988E+03    4

HNO2                    H   1N   1O   2     G  0300.00   4000.00  1500.00      1 ! RASMUSSEN 2008; Int J Chem Kinet 40: 454â€“480, 2008(ab initio CBS-QB3); 

 6.47963000E+00 1.99527400E-03-1.74038700E-07-9.69587200E-11 1.70148000E-14    2 ! H298=-9.80 kcal/mol

-7.80950291E+03-1.06771518E+01 1.93483800E+00 1.01003600E-02-4.96461600E-06    3 ! S298=56.73 cal/mol/K [Sandia]

 8.70112000E-10-2.32413500E-15-5.91571591E+03 1.47282082E+01                   4 !

HONO2             T 8/03H   1N   1O   3    0G   200.00   6000.00  1000.        1 ! RASMUSSEN 2008; Int J Chem Kinet 40: 454â€“480, 2008

 8.03098942E+00 4.46958589E-03-1.72459491E-06 2.91556153E-10-1.80102702E-14    2 ! H298 = -134.112+/-0.18 kJ/mol 

-1.92821685E+04-1.62616720E+01 1.69329154E+00 1.90167702E-02-8.25176697E-06    3 ! S298 = 63.76 cal/mol/K 

-6.06113827E-09 4.65236978E-12-1.73882411E+04 1.71839655E+01                   4 

NO3               ATcT/AN   1O   3    0    0G   200.00   6000.00  1000.0       1 ! Burcat/Goos 2017

 7.48347702E+00 2.57772064E-03-1.00945831E-06 1.72314063E-10-1.07154008E-14    2 

 6.12990474E+03-1.41618136E+01 2.17359330E+00 1.04902685E-02 1.10472669E-05    3 

-2.81561867E-08 1.36583960E-11 7.81290905E+03 1.46022090E+01 8.97563416E+03    4 

N2O3              L 4/90N   2O   3    0    0G   200.000  6000.000 1000.        1 ! Burcat/Goos 2017

 9.08583845E+00 3.37756330E-03-1.31583890E-06 2.30762329E-10-1.47151267E-14    2

 7.27160146E+03-1.55361904E+01 5.81083964E+00 1.43330962E-02-1.96208597E-05    3

 1.73060735E-08-6.46553954E-12 8.19184453E+03 1.20461321E+00 1.04192062E+04    4

N2O4              ATcT AN  2.O  4.   0.   0.G   200.000  6000.000 1000.        1 ! Burcat/Goos 2017

 1.15752932E+01 4.01615532E-03-1.57178022E-06 2.68273657E-10-1.66921538E-14    2

-2.96111235E+03-3.19488625E+01 3.02002271E+00 2.95904359E-02-3.01342572E-05    3

 1.42360526E-08-2.44100411E-12-6.79238803E+02 1.18059620E+01 1.29712996E+03    4 

HNO3              T 8/03H  1.N  1.O  3.   0.G   200.000  6000.000 1000.        1 ! Burcat/Goos 2017

 8.03098942E+00 4.46958589E-03-1.72459491E-06 2.91556153E-10-1.80102702E-14    2

-1.93138183E+04-1.62616537E+01 1.69329154E+00 1.90167702E-02-8.25176697E-06    3

-6.06113827E-09 4.65236978E-12-1.74198909E+04 1.71839838E+01-1.61524852E+04    4

CH3ONO            A 5/05C   1H   3O   2N   1G   200.00   6000.00  1000.0       1 ! Burcat/Goos 2017 ! Methyl-Nitrite

 6.93605239E+00 9.97319424E-03-3.60642537E-06 5.83462161E-10-3.50058729E-14    2

-1.08381899E+04-6.98144573E+00 6.15261387E+00-2.91937431E-03 4.14526828E-05    3

-4.93954776E-08 1.85608328E-11-9.85260262E+03 8.04057190E-01-7.87057806E+03    4

CH3NO NitrosomethyT12/09C  1.H  3.N  1.O  1.G   200.000  6000.000 1000.0       1 ! Burcat/Goos 2017 ! NITROSOMETHYL or METHYL-NITROSYL

 5.04711802E+00 9.21544305E-03-3.29034831E-06 5.28940397E-10-3.15689858E-14    2

 6.23718102E+03-7.74395570E-01 5.18534727E+00-6.34085575E-03 4.57171139E-05    3

-5.30421813E-08 1.99501601E-11 6.93771506E+03 2.18492659E+00 8.51040025E+03    4

CH3ONO2           T05/98C   1H   3N   1O   3G   200.00   6000.00  1000.0       1 ! Burcat/Goos 2017 ! Methyl-Nitrate

 9.77845489E+00 1.10069541E-02-4.25928645E-06 7.18198185E-10-4.42041793E-14    2 

-1.88804487E+04-2.39163197E+01 3.91363583E+00 1.52137945E-02 1.73479131E-05    3 

-3.37074473E-08 1.44322204E-11-1.66103232E+04 9.44208392E+00-1.46737980E+04    4

CH3NO2            T01/00C   1H   3N   1O   2G   200.000  6000.000 1000.0       1 ! Burcat/Goos 2017 ! Nitro-Methane

 6.73034758E+00 1.09601272E-02-4.05357875E-06 6.67102246E-10-4.04686823E-14    2

-1.29143475E+04-1.01800883E+01 3.54053638E+00 1.86559899E-03 4.44946580E-05    3

-5.87057133E-08 2.30684496E-11-1.11385976E+04 1.06884657E+01-9.71208165E+03    4

CH2NO2  RADICAL  T08/07 C  1.H  2.N  1.O  2.G   200.000  6000.000 1000.0       1 ! Burcat/Goos 2017

 7.57504807E+00 7.01471036E-03-2.51481162E-06 4.05670550E-10-2.42796598E-14    2

 1.23880080E+04-1.15985589E+01 2.42742248E+00 1.60496442E-02 2.84727836E-06    3

-1.82218429E-08 9.35383557E-12 1.40120587E+04 1.61086425E+01 1.54427130E+04    4

CH2CN   BUR0302   T01/03C  2.H  2.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat/Goos 2017

 6.14873620E+00 6.06600240E-03-2.17174620E-06 3.49750387E-10-2.09004207E-14    2 ! METHYLENECYANIDE RADICAL

 2.86491222E+04-6.59235995E+00 2.63064017E+00 1.73644377E-02-1.70284117E-05    3

 9.86551140E-09-2.46033517E-12 2.95791691E+04 1.12776223E+01 3.10031788E+04    4

CH3CN  BUR0302    T01/03C  2.H  3.N  1.   0.G   200.000  6000.000 1000.        1 ! Burcat/Goos 2017

 5.09921882E+00 9.69585649E-03-3.48051966E-06 5.61420173E-10-3.35835856E-14    2 ! METHYLCYANIDE 

 6.60967324E+03-3.36087178E+00 3.82392803E+00 4.08201943E-03 2.16209537E-05    3 !

-2.89807789E-08 1.12962700E-11 7.44430382E+03 5.52656156E+00 8.90492212E+03    4

!CH2NO  H2C=N-O*   T06/08C  1.H  2.N  1.O  1.G   200.000  6000.000 1000.        1 ! Burcat 2017

! 5.41478025E+00 6.68230119E-03-2.38625695E-06 3.83764001E-10-2.29149657E-14    2

! 1.63459530E+04-3.03719498E+00 3.00389272E+00 6.88209471E-03 1.26563213E-05    3

!-2.17579528E-08 9.28731765E-12 1.73161337E+04 1.09485576E+01 1.85908365E+04    4

!CH2NO H2C*N=O RADICAL The G3B3 calculations show that this conformation is in   !

!resonance with the former conformation H2C*N=O <=> H2C=M-O* therefore the former!

!polynomial should be used here. The present polynomial comes from the data of   !

!C. Melius BAC/MP4 calculations of 1987.  STATWT=2  SIGMA=2  IA=2.596  IB=3.041  !

!IC=5.0754   NU=3040,2952,1505,1304,1188,1111,983,897,846   HF298=53.52+/-2 kcal !

!REF=C. MELIUS DATABASE BAC/MP4 D93X  Max Lst Sq Error Cp @ 200 K 0.82%.

CH2NO  H2C*N=O    T 9/96C   1H   2N   1O   1G    200.00   6000.00 1000.00      1 ! E. Goos, A. Burcat, and B. Ruscic

 0.54028152E+01 0.69057001E-02-0.25162977E-05 0.41014066E-09-0.24718300E-13    2 ! Ideal gas thermochemical database with updates from active thermochemical

 0.24528690E+05-0.44574262E+01 0.38781858E+01-0.66530886E-02 0.53947610E-04    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

-0.68176813E-07 0.27181746E-10 0.25716857E+05 0.74618774E+01 0.26932156E+05    4 ! Accessed 2018

!CH2NO       MELIUS 88   H   2N   1C   1O   1G   300.000  5000.000 1394.000     1 ! He 2016

! 6.93551152E+00 5.19106959E-03-1.80090529E-06 2.82284906E-10-1.64876420E-14    2 

! 1.78889823E+04-1.16990566E+01 1.35048335E+00 1.95270193E-02-1.62924222E-05    3 

! 7.08039958E-09-1.24896699E-12 1.97105070E+04 1.78571822E+01                   4 

HON          HF MELIUS93H   1N   1O   1    0G   300.000  5000.000 1671.000     1 ! Mathieu et al 2016; Fuel 182 (2016) 597â€“612

 3.78577430E+00 2.86062728E-03-1.02423922E-06 1.64463139E-10-9.77943616E-15    2

 2.93319701E+04 3.12193293E+00 3.33656431E+00 2.67682939E-03 5.61801303E-07    3

-1.11362279E-09 2.84076438E-13 2.95979751E+04 5.96343188E+00                   4

!HON                     H   1N   1O   1     G   298.150  3000.000 1000.00      1 ! Bugler 2016; J. Phys. Chem. A 2016, 120, 7192âˆ’7197

! 3.71174626E+00 3.16088951E-03-1.33270405E-06 2.82287945E-10-2.37381901E-14    2

! 2.44108221E+04 5.58114551E+00 3.05581786E+00 4.43591111E-03-1.22219840E-06    3

!-1.14007451E-09 6.69025432E-13 2.46094424E+04 9.08279393E+00                   4

!CH3NH2      SWS         H   5C   1N   1    0G   300.000  5000.000 1387.000     1 ! DB00

! 5.23365618E+00 1.08525479E-02-3.65205276E-06 5.60552543E-10-3.22553444E-14    2 ! Mathieu et al. 2016; Fuel 182 (2016) 597â€“612

!-5.52829576E+03-5.21507359E+00 1.69170293E+00 1.60389160E-02-4.99028441E-06    3

!-3.83481304E-10 3.57345746E-13-3.94057426E+03 1.49835076E+01                   4

CH3NH2            T09/09C  1.H  5.N  1.   0.G   200.000  6000.000 1000.        1 ! METHYLAMINE ! E. Goos, A. Burcat, and B. Ruscic

 3.78609899E+00 1.26969570E-02-4.46778553E-06 7.11021516E-10-4.21332621E-14    2 ! Ideal gas thermochemical database with updates from active thermochemical

-4.38100060E+03 1.86268606E+00 4.65718252E+00-7.37953092E-03 5.45297099E-05    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

-6.24993857E-08 2.33761829E-11-3.76073340E+03 1.63875112E+00-2.33089960E+03    4 ! Accessed 2018

!CH3NH       THERM92     H   4C   1N   1    0G   300.000  5000.000 1404.000     1 ! DB00

! 4.90528413E+00 8.50385569E-03-2.82356461E-06 4.29267836E-10-2.45297886E-14    2 ! Mathieu et al. 2016; Fuel 182 (2016) 597â€“612

! 1.94541503E+04-1.35290137E+00 1.53882571E+00 1.62436539E-02-9.89573425E-06    3

! 3.49954504E-09-5.53823621E-13 2.06715086E+04 1.68295527E+01                   4

CH3NH radical     T03/10C  1.H  4.N  1.   0.G   200.000  6000.000 1000.        1 ! METHYL AMINO RADICAL ! E. Goos, A. Burcat, and B. Ruscic

 4.02244380E+00 1.03512061E-02-3.64560169E-06 5.80491587E-10-3.44103829E-14    2 ! Ideal gas thermochemical database with updates from active thermochemical

 1.95050854E+04 1.64483768E+00 4.70973738E+00-7.31946952E-03 4.95105509E-05    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

-5.72790480E-08 2.16523586E-11 2.00619432E+04 1.85460205E+00 2.14752744E+04    4 ! Accessed 2018

!CH2NH2      THERM92     H   4C   1N   1    0G   300.000  5000.000 1397.000     1 ! DB00

! 6.11432288E+00 7.69126269E-03-2.59025729E-06 3.97713575E-10-2.28883272E-14    2 ! Mathieu et al. 2016; Fuel 182 (2016) 597â€“612

! 1.55835138E+04-8.93053780E+00 2.56157769E+00 1.60730713E-02-1.05960335E-05    3 ! He et al. 2016; Energy Fuels 2016, 30, 6799âˆ’6807

! 4.07638829E-09-6.95570548E-13 1.68563722E+04 1.01987687E+01                   4

CH2NH2 radical    T03/10C   1H   4N  1     0G    200.00  6000.00 1000.0        1 ! MethenyAmine AminoMethyl Radical; E. Goos, A. Burcat, and B. Ruscic

 4.55329728E+00 9.42002581E-03-3.20781399E-06 4.98961894E-10-2.90872284E-14    2 ! Ideal gas thermochemical database with updates from active thermochemical

 1.58717284E+04-2.45945234E-02 2.85538164E+00 7.27364238E-03 1.65712636E-05    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

-2.70976978E-08 1.16327939E-11 1.66165986E+04 1.02444521E+01 1.78895690E+04    4 ! Accessed 2018

!CH2NH       MELIUS 88   H   3C   1N   1    0G   300.000  5000.000 1577.000     1 ! DB00

! 4.54737795E+00 7.17720948E-03-2.47935299E-06 3.87692351E-10-2.26113075E-14    2 ! Mathieu et al. 2016; Fuel 182 (2016) 597â€“612

! 8.64056516E+03-1.16687427E+00 2.81849510E+00 5.11983235E-03 6.38887146E-06    3

!-6.61374671E-09 1.65531940E-12 9.88442597E+03 1.03390629E+01                   4

CH2NH  (H2C=NH)   A12/04H   3C   1N   1    0G   200.000  6000.000 1000.        1 ! METHANIMINE ! E. Goos, A. Burcat, and B. Ruscic

 3.44258358E+00 8.37600036E-03-2.97819078E-06 4.77352867E-10-2.84295062E-14    2 ! Ideal gas thermochemical database with updates from active thermochemical

 8.40771949E+03 3.95595397E+00 4.79302577E+00-1.26841692E-02 5.69766521E-05    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

-6.34985251E-08 2.37023330E-11 8.85023146E+03 1.10277996E+00 1.01045906E+04    4 ! Accessed 2018 

!HCNH               41687C   1H   2N   1     G  0300.00   4000.00  1000.00      1 ! Mathieu et al. 2016; Fuel 182 (2016) 597â€“612

! 0.04923293E+02 0.03332897E-01-0.03370897E-05-0.01901619E-08 0.03531825E-12    2

! 0.03132669E+06-0.01632509E+02 0.02759456E+02 0.06103387E-01 0.07713149E-05    3

!-0.02063094E-07 0.01931920E-11 0.03217247E+06 0.01057489E+03                   4

HCNH  H*C=NH Tra  T10/09C  1.H  2.N  1.   0.G   200.000  6000.000 1000.        1 ! (H*C=NH) RADICAL trans; ! E. Goos, A. Burcat, and B. Ruscic

 4.04014700E+00 5.16591694E-03-1.82276828E-06 2.90299053E-10-1.71614589E-14    2 ! Ideal gas thermochemical database with updates from active thermochemical

 3.42988367E+04 2.58894095E+00 3.97114555E+00-3.88875724E-03 2.92918950E-05    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

-3.57482411E-08 1.40303911E-11 3.47237453E+04 5.06388721E+00 3.59296699E+04    4 ! Accessed 2018 

! It is strictly forbidden to include this database as it is or parts of it    !

! in any commercial database, software, firmware or hardware and any other type!

! of commercial use without written permission from the authors. For commercial!

! use and non combustion relevant substances please contact info@thermodata.de !

!HCNH  H*C=NH  cis T10/09C  1.H  2.N  1.   0.G   200.000  6000.000 1000.        1 ! (H*C=NH) RADICAL cis; ! E. Goos, A. Burcat, and B. Ruscic

! 4.21964637E+00 5.00385318E-03-1.76392242E-06 2.80726369E-10-1.65852271E-14    2 ! Ideal gas thermochemical database with updates from active thermochemical

! 3.67706425E+04 1.67137973E+00 3.68324272E+00-1.38553491E-03 2.40042193E-05    3 ! http://garfield.chem.elte.hu/Burcat/burcat.html

!-3.11573911E-08 1.25791822E-11 3.72527355E+04 6.21247271E+00 3.84457533E+04    4 ! Accessed 2018 





! Thermo (not BAC corrected because I do not have those for nitrogen compounds)

!        (could develop those if needed)   

! {SpName = IPN }  { IPN }

! {3Freq =   362.257  11.672  1196.232  15.569  2708.376   6.759  }

! {LJepsilon = xxx }  {LJsigma = xxx }  {KMOI = 1.23 }

! {E0 =   -43.14 }  {CalcMeth = CBS-QB3 }                                                                                                 

IPN               092619H   7C   3N   1O   3g   300.000  2500.000 1000.000     1

 0.71500983E+01 0.39662939E-01-0.22521714E-04 0.62039458E-08-0.67388358E-12    2

-0.29119332E+05-0.78215566E+01 0.16013503E+01 0.50701205E-01-0.20059560E-04    3

-0.10562923E-07 0.81436299E-11-0.27482219E+05 0.21623074E+02           HHC 4 P 4

 

! {SpName = CH2CHCH3ONO2 }  { CH2CHCH3ONO2 }

! {3Freq =   361.255  12.570  1243.787  13.437  2905.347   4.993  }

! {LJepsilon = xxx }  {LJsigma = xxx }  {KMOI = 1.23 }

! {E0 =     6.90 }  {CalcMeth = CBS-QB3 } 

CH2CHCH3ONO2      042220H   6C   3N   1O   3g   300.000  2500.0001000.000      1

 0.91725359E+01 0.32913681E-01-0.18622341E-04 0.51259423E-08-0.55716488E-12    2

-0.35658865E+04-0.14982266E+02 0.28678088E+01 0.48613671E-01-0.26154430E-04    3

-0.24695492E-08 0.51770892E-11-0.18484358E+04 0.17733568E+02           HHC 4 M 4

CH3CHOCH2               C   3H   6O   1     G  0300.00   5000.00  1000.00      1

 0.91590881E+01 0.15399657E-01-0.51697507E-05 0.81830304E-09-0.50199259E-13    2

-0.15840833E+05-0.24935184E+02 0.77822632E+00 0.29787362E-01-0.11344674E-04    3

 0.86544716E-09 0.63418163E-13-0.12630026E+05 0.21613398E+02                   4

IC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1527.000    21

 1.19648494E+01 1.42943974E-02-4.71413211E-06 7.14027066E-10-4.07161162E-14    2

-1.17519389E+04-3.88860959E+01 2.36108410E+00 3.45650027E-02-1.94579631E-05    3

 4.71536901E-09-2.64704937E-13-8.28791395E+03 1.33112436E+01                   4

CH3COCH3   8/12/15      C   3H   6O   1    0G   300.000  5000.000 1394.000    21

 8.87619308E+00 1.45700263E-02-4.84823280E-06 7.38614777E-10-4.22831194E-14    2

-3.06046242E+04-2.12730484E+01 2.20008426E+00 2.74019559E-02-1.31342003E-05    3

 2.57150371E-09-6.21509091E-14-2.79933966E+04 1.55883508E+01                   4

IC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1000.00      1

 .964183701E+01 .200230715E-01-.711967189E-05 .114138950E-08-.679935249E-13    2

-.374835623E+05-.256288343E+02 .430755345E+01 .102582798E-01 .619565411E-04    3

-.902973802E-07 .373936384E-10-.349249212E+05 .755995822E+01                   4

CH3COCH2   2/14/13 THERMC   3H   5O   1    0G   300.000  5000.000 1387.000    21

 1.09524298E+01 1.11458668E-02-3.86262877E-06 6.05088857E-10-3.53293362E-14    2

-9.60833727E+03-3.15622776E+01 1.13381826E+00 3.25095045E-02-2.10424651E-05    3

 6.64421151E-09-8.12618901E-13-6.04868361E+03 2.17158655E+01                   4

HOCO       9/27/ 5 THERMC   1H   1O   2    0G   300.000  5000.000 1549.000    11

 6.94282268E+00 2.37391844E-03-8.67074662E-07 1.40644617E-10-8.41268695E-15    2

-2.50292163E+04-1.14792361E+01 8.98154532E-01 1.67269019E-02-1.33663562E-05    3

 4.83071199E-09-6.38718748E-13-2.30262021E+04 2.07803865E+01                   4



END



















