!VERSION:  16_03
!AUTHORS:  C3
!NOTE:     SPECIES RE-ARRANGED AS THE SAME ORDER IN MECH
THERMO
   300.000  1000.000  5000.000
AR                G 5/97AR  1  0    0      0G   200.000  6000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 4.37967491E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 4.37967491E+00 0.00000000E+00    4
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
HE                G 5/97HE 1    0    0    0 G   200.000  6000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 9.28723974E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 9.28723974E-01 0.00000000E+00    4
H2                TPIS78H   2    0    0    0G   200.000  6000.00  1000.00      1
 2.93286575E+00 8.26608026E-04-1.46402364E-07 1.54100414E-11-6.88804800E-16    2
-8.13065581E+02-1.02432865E+00 2.34433112E+00 7.98052075E-03-1.94781510E-05    3
 2.01572094E-08-7.37611761E-12-9.17935173E+02 6.83010238E-01 0.00000000E+00    4
H                 L 6/94H   1    0    0    0G   200.000  6000.00  1000.00      1
 0.25000000E+01 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.25473660E+05-0.44668285E+00 0.25000000E+01 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.25473660E+05-0.44668285E+00 0.26219035E+05    4
O2                RUS 89O   2    0    0    0G   200.000  6000.00  1000.00      1
 3.66096065E+00 6.56365811E-04-1.41149627E-07 2.05797935E-11-1.29913436E-15    2
-1.21597718E+03 3.41536279E+00 3.78245636E+00-2.99673416E-03 9.84730201E-06    3
-9.68129509E-09 3.24372837E-12-1.06394356E+03 3.65767573E+00 0.00000000E+00    4
O                 L 1/90O   1    0    0    0G   200.000  6000.00  1000.00      1
 2.54363697E+00-2.73162486E-05-4.19029520E-09 4.95481845E-12-4.79553694E-16    2
 2.92260120E+04 4.92229457E+00 3.16826710E+00-3.27931884E-03 6.64306396E-06    3
-6.12806624E-09 2.11265971E-12 2.91222592E+04 2.05193346E+00 2.99687009E+04    4
H2O               L 5/89H   2 O  1    0    0G   200.000  6000.00  1000.00      1
 0.26770389E+01 0.29731816E-02-0.77376889E-06 0.94433514E-10-0.42689991E-14    2
-0.29885894E+05 0.68825500E+01 0.41986352E+01-0.20364017E-02 0.65203416E-05    3
-0.54879269E-08 0.17719680E-11-0.30293726E+05-0.84900901E+00-0.29084817E+05    4
OH                IU3/03O   1 H  1    0    0G   200.000  6000.00  1000.00      1
 2.83853033E+00 1.10741289E-03-2.94000209E-07 4.20698729E-11-2.42289890E-15    2
 3.69780808E+03 5.84494652E+00 3.99198424E+00-2.40106655E-03 4.61664033E-06    3
-3.87916306E-09 1.36319502E-12 3.36889836E+03-1.03998477E-01 4.48613328E+03    4
OHV               121286O   1H   1          G  0300.00   5000.00  1000.00      1
 0.02882730E+02 0.10139743E-02-0.02276877E-05 0.02174683E-09-0.05126305E-14    2
 5.02650000E+04 0.05595712E+02 0.03637266E+02 0.01850910E-02-0.16761646E-05    3
 0.02387202E-07-0.08431442E-11 5.00213000E+04 0.13588605E+01                   4
H2O2              T 8/03H   2O   2    0    0G   200.000  6000.00  1000.00      1
 4.57977305E+00 4.05326003E-03-1.29844730E-06 1.98211400E-10-1.13968792E-14    2
-1.80071775E+04 6.64970694E-01 4.31515149E+00-8.47390622E-04 1.76404323E-05    3
-2.26762944E-08 9.08950158E-12-1.77067437E+04 3.27373319E+00-1.63425145E+04    4
HO2               T 1/09H   1O   2    0    0G   200.000  5000.00  1000.00      1
 4.17228741E+00 1.88117627E-03-3.46277286E-07 1.94657549E-11 1.76256905E-16    2
 3.10206839E+01 2.95767672E+00 4.30179807E+00-4.74912097E-03 2.11582905E-05    3
-2.42763914E-08 9.29225225E-12 2.64018485E+02 3.71666220E+00 1.47886045E+03    4
CO                RUS 79C   1O   1    0    0G   200.000  6000.00  1000.00      1
 0.30484859E+01 0.13517281E-02-0.48579405E-06 0.78853644E-10-0.46980746E-14    2
-0.14266117E+05 0.60170977E+01 0.35795335E+01-0.61035369E-03 0.10168143E-05    3
 0.90700586E-09-0.90442449E-12-0.14344086E+05 0.35084093E+01-0.13293628E+05    4
CO2               L 7/88C   1O   2    0    0G   200.000  6000.00  1000.00      1
 0.46365111E+01 0.27414569E-02-0.99589759E-06 0.16038666E-09-0.91619857E-14    2
-0.49024904E+05-0.19348955E+01 0.23568130E+01 0.89841299E-02-0.71220632E-05    3
 0.24573008E-08-0.14288548E-12-0.48371971E+05 0.99009035E+01-0.47328105E+05    4
HOCO              T05/06H  1 C  1 O  2    0 G   200.000  6000.00   1000.00     1
 5.39206152E+00 4.11221455E-03-1.48194900E-06 2.39875460E-10-1.43903104E-14    2
-2.38606717E+04-2.23529091E+00 2.92207919E+00 7.62453859E-03 3.29884437E-06    3
-1.07135205E-08 5.11587057E-12-2.30281524E+04 1.12925886E+01-2.18076591E+04    4
CH4               G 8/99C  1 H  4    0    0 G   200.000  6000.00  1000.00      1
 1.65326226E+00 1.00263099E-02-3.31661238E-06 5.36483138E-10-3.14696758E-14    2
-1.00095936E+04 9.90506283E+00 5.14911468E+00-1.36622009E-02 4.91453921E-05    3
-4.84246767E-08 1.66603441E-11-1.02465983E+04-4.63848842E+00-8.97226656E+03    4
CH3               IU0702C  1 H  3    0    0 G   200.000  6000.00  1000.00      1
 0.29781206E+01 0.57978520E-02-0.19755800E-05 0.30729790E-09-0.17917416E-13    2
 0.16509513E+05 0.47224799E+01 0.36571797E+01 0.21265979E-02 0.54583883E-05    3
-0.66181003E-08 0.24657074E-11 0.16422716E+05 0.16735354E+01 0.17643935E+05    4
CH2               IU3/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
 3.14631886E+00 3.03671259E-03-9.96474439E-07 1.50483580E-10-8.57335515E-15    2
 4.60412605E+04 4.72341711E+00 3.71757846E+00 1.27391260E-03 2.17347251E-06    3
-3.48858500E-09 1.65208866E-12 4.58723866E+04 1.75297945E+00 4.70504920E+04    4
CH2(S)            IU6/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
 3.13501686E+00 2.89593926E-03-8.16668090E-07 1.13572697E-10-6.36262835E-15    2
 5.05040504E+04 4.06030621E+00 4.19331325E+00-2.33105184E-03 8.15676451E-06    3
-6.62985981E-09 1.93233199E-12 5.03662246E+04-7.46734310E-01 5.15727280E+04    4
C                 L 7/88C   1     0    0   0G   200.000  6000.00  1000.00      1
 0.26055830E+01-0.19593434E-03 0.10673722E-06-0.16423940E-10 0.81870580E-15    2
 0.85411742E+05 0.41923868E+01 0.25542395E+01-0.32153772E-03 0.73379223E-06    3
-0.73223487E-09 0.26652144E-12 0.85442681E+05 0.45313085E+01 0.86195097E+05    4
CH                IU3/03C  1 H  1    0    0 G   200.000  6000.00  1000.00      1
 0.25209369E+01 0.17653639E-02-0.46147660E-06 0.59289675E-10-0.33474501E-14    2
 0.70946769E+05 0.74051829E+01 0.34897583E+01 0.32432160E-03-0.16899751E-05    3
 0.31628420E-08-0.14061803E-11 0.70612646E+05 0.20842841E+01 0.71658188E+05    4
CHV               073003C   1H   1          G  0300.00   5000.00  1000.00      1
 0.02196223E+02 0.02340381E-01-0.07058201E-05 0.09007582E-09-0.03855040E-13    2
 0.10419559E+06 0.09178373E+02 0.03200202E+02 0.02072875E-01-0.05134431E-04    3
 0.05733890E-07-0.01955533E-10 0.10393714E+06 0.03331587E+02                   4
CH3O2H            A 7/05C  1 H  4 O  2    0 G   200.000  6000.00  1000.00      1
 7.76538058E+00 8.61499712E-03-2.98006935E-06 4.68638071E-10-2.75339255E-14    2
-1.82979984E+04-1.43992663E+01 2.90540897E+00 1.74994735E-02 5.28243630E-06    3
-2.52827275E-08 1.34368212E-11-1.68894632E+04 1.13741987E+01-1.52423685E+04    4
CH3O2                   H   3C   1O   2    0G   300.000  5000.000 1374.000     1
 6.47970487E+00 7.44401080E-03-2.52348555E-06 3.89577296E-10-2.25182399E-14    2
-1.56285441E+03-8.19477074E+00 1.97339205E+00 1.53542340E-02-6.37314891E-06    3
 3.19930565E-10 2.82193915E-13 2.54278835E+02 1.69194215E+01                   4
CH2O2H     9/ 1/12      C   1H   3O   2    0G   300.000  5000.000 1410.000     1
 9.24697852E+00 4.60845541E-03-1.53501472E-06 2.34434830E-10-1.34573106E-14    2
 4.11529953E+03-2.11503248E+01 2.88976454E+00 2.09465776E-02-1.75190772E-05    3
 7.27819787E-09-1.18912344E-12 6.12390620E+03 1.23802076E+01                   4
CH3OH             T06/02C   1H  4 O  1    0 G   200.000  6000.00  1000.00      1
 3.52726795E+00 1.03178783E-02-3.62892944E-06 5.77448016E-10-3.42182632E-14    2
-2.60028834E+04 5.16758693E+00 5.65851051E+00-1.62983419E-02 6.91938156E-05    3
-7.58372926E-08 2.80427550E-11-2.56119736E+04-8.97330508E-01-2.41746056E+04    4
CH3O              IU1/03C  1 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 4.75779238E+00 7.44142474E-03-2.69705176E-06 4.38090504E-10-2.63537098E-14    2
 3.78111940E+02-1.96680028E+00 3.71180502E+00-2.80463306E-03 3.76550971E-05    3
-4.73072089E-08 1.86588420E-11 1.29569760E+03 6.57240864E+00 2.52571660E+03    4
CH2OH             IU2/03C  1 H  3 O  1    0 G   200.000  6000.00   1000.00     1
 5.09314370E+00 5.94761260E-03-2.06497460E-06 3.23008173E-10-1.88125902E-14    2
-4.03409640E+03-1.84691493E+00 4.47834367E+00-1.35070310E-03 2.78484980E-05    3
-3.64869060E-08 1.47907450E-11-3.50072890E+03 3.30913500E+00-2.04462770E+03    4
CH2O              T 5/11H   2C   1O   1    0G   200.000  6000.00  1000.00      1
 3.16952665E+00 6.19320560E-03-2.25056366E-06 3.65975660E-10-2.20149458E-14    2
-1.45486831E+04 6.04207898E+00 4.79372312E+00-9.90833322E-03 3.73219990E-05    3
-3.79285237E-08 1.31772641E-11-1.43791953E+04 6.02798058E-01-1.31293365E+04    4
HCO               T 5/03C  1 H  1 O  1    0 G   200.000  6000.00  1000.00      1
 3.92001542E+00 2.52279324E-03-6.71004164E-07 1.05615948E-10-7.43798261E-15    2
 3.65342928E+03 3.58077056E+00 4.23754610E+00-3.32075257E-03 1.40030264E-05    3
-1.34239995E-08 4.37416208E-12 3.87241185E+03 3.30834869E+00 5.08749163E+03    4
HCOH              MAR94 C   1H   2O   1    0G   300.     5000.    1398.        1
 9.18749272E+00 1.52011152E-03-6.27603516E-07 1.09727989E-10-6.89655128E-15    2
 7.81364593E+03-2.73434214E+01-2.82157421E+00 3.57331702E-02-3.80861580E-05    3
 1.86205951E-08-3.45957838E-12 1.12956672E+04 3.48487757E+01                   4
HO2CHO     6/26/95 THERMC   1H   2O   3    0G   300.000  5000.000 1378.00      1
 9.87503878E+00 4.64663708E-03-1.67230522E-06 2.68624413E-10-1.59595232E-14    2
-3.80502496E+04-2.24939155E+01 2.42464726E+00 2.19706380E-02-1.68705546E-05    3
 6.25612194E-09-9.11645843E-13-3.54828006E+04 1.75027796E+01                   4
HOCH2O2H   9/ 1/12      C   1H   4O   3    0G   300.000  5000.000 1398.000     1
 1.24531886E+01 7.18221110E-03-2.47029548E-06 3.85611737E-10-2.24774193E-14    2
-4.24862928E+04-3.58745197E+01 5.35189713E-01 3.73266553E-02-3.15299511E-05    3
 1.30352583E-08-2.11473264E-12-3.86609415E+04 2.71776082E+01                   4
HOCH2O2    9/ 1/12      C   1H   3O   3    0G   300.000  5000.000 1377.000     1
 1.16406115E+01 5.72826040E-03-2.05362036E-06 3.29070695E-10-1.95188360E-14    2
-2.53505769E+04-3.07332064E+01 2.82068616E+00 2.47857094E-02-1.66186399E-05    3
 4.79633095E-09-4.28087766E-13-2.22077036E+04 1.70599803E+01                   4
OCH2O2H    7/21/14 THERMC   1H   3O   3    0G   300.000  5000.000 1418.000     1
 1.29622491E+01 4.21948855E-03-1.54275194E-06 2.50413077E-10-1.49855537E-14    2
-1.81326406E+04-3.87016356E+01 4.46349361E-01 3.63049606E-02-3.26130978E-05    3
 1.37050551E-08-2.20872791E-12-1.41972598E+04 2.72960376E+01                   4
HOCH2O     2/16/99 THERMC   1H   3O   2    0G   300.000  5000.000 1452.000     1
 6.39521515E+00 7.43673043E-03-2.50422354E-06 3.84879712E-10-2.21778689E-14    2
-2.41108840E+04-6.63865583E+00 4.11183145E+00 7.53850697E-03 3.77337370E-06    3
-5.38746005E-09 1.45615887E-12-2.28023001E+04 7.46807254E+00                   4
O2CHO      6/26/95 THERMC   1H   1O   3    0G   300.000  5000.000 1368.00      1
 7.24075139E+00 4.63312951E-03-1.63693995E-06 2.59706693E-10-1.52964699E-14    2
-1.87027618E+04-6.49547212E+00 3.96059309E+00 1.06002279E-02-5.25713351E-06    3
 1.01716726E-09-2.87487602E-14-1.73599383E+04 1.17807483E+01                   4
HOCHO             L 8/88H   2C   1O   2    0G   200.000  6000.00  1000.00      1
 0.46138316E+01 0.64496364E-02-0.22908251E-05 0.36716047E-09-0.21873675E-13    2
-0.47514850E+05 0.84788383E+00 0.38983616E+01-0.35587795E-02 0.35520538E-04    3
-0.43849959E-07 0.17107769E-10-0.46770609E+05 0.73495397E+01-0.45531246E+05    4
OCHO              ATCT/AC  1 O  2 H  1    0 G   200.000  6000.000 1000.00      1
 4.14394211E+00 5.59738818E-03-1.99794019E-06 3.16179193E-10-1.85614483E-14    2
-1.72459887E+04 5.07778617E+00 4.68825921E+00-4.14871834E-03 2.55066010E-05    3
-2.84473900E-08 1.04422559E-11-1.69867041E+04 4.28426480E+00-1.55992356E+04    4
C2H6              G 8/88C   2H 6    0      0G   200.000  6000.00  1000.00      1
 4.04666411E+00 1.53538802E-02-5.47039485E-06 8.77826544E-10-5.23167531E-14    2
-1.24473499E+04-9.68698313E-01 4.29142572E+00-5.50154901E-03 5.99438458E-05    3
-7.08466469E-08 2.68685836E-11-1.15222056E+04 2.66678994E+00-1.00849652E+04    4
C2H5       8/ 4/ 4 THERMC   2H   5    0    0G   300.000  5000.000 1387.000     1
 5.88784390E+00 1.03076793E-02-3.46844396E-06 5.32499257E-10-3.06512651E-14    2
 1.15065499E+04-8.49651771E+00 1.32730217E+00 1.76656753E-02-6.14926558E-06    3
-3.01143466E-10 4.38617775E-13 1.34284028E+04 1.71789216E+01                   4
C2H5O2H    9/ 1/12      C   2H   6O   2    0G   300.000  5000.000 1390.000     1
 1.04823538E+01 1.34779879E-02-4.62179078E-06 7.18618519E-10-4.17307436E-14    2
-2.46578171E+04-2.84294243E+01 1.83755328E+00 3.38053586E-02-2.37548140E-05    3
 9.31974865E-09-1.58003428E-12-2.15814086E+04 1.80977584E+01                   4
C2H5O2     9/ 1/12      C   2H   5O   2    0G   300.000  5000.000 1389.000     1
 9.50282570E+00 1.20429839E-02-4.09491581E-06 6.33049241E-10-3.66133788E-14    2
-7.37069391E+03-2.21717130E+01 3.90351912E+00 2.22599212E-02-1.01610079E-05    3
 1.71709751E-09 1.88166738E-14-5.09654081E+03 8.98722750E+00                   4
C2H4       8/12/15      C   2H   4    0    0G   300.000  5000.000 1392.000     1
 5.07061289E+00 9.11140768E-03-3.10506692E-06 4.80733851E-10-2.78321396E-14    2
 3.66391217E+03-6.64501414E+00 4.81118223E-01 1.83778060E-02-9.99633565E-06    3
 2.73211039E-09-3.01837289E-13 5.44386648E+03 1.85867157E+01                   4
C2H3       8/12/15      C   2H   3    0    0G   300.000  5000.000 1400.000     1
 4.99675415E+00 6.55838271E-03-2.20921909E-06 3.39300272E-10-1.95316926E-14    2
 3.34604382E+04-3.01451097E+00 1.25545094E+00 1.57481597E-02-1.12218328E-05    3
 4.50915682E-09-7.74861577E-13 3.47435574E+04 1.69664043E+01                   4
CHOCHO                  C   2H   2O   2    0G   300.000  5000.000 1386.000     1
 9.75438561E+00 4.97645947E-03-1.74410483E-06 2.75586994E-10-1.61969892E-14    2
-2.95832896E+04-2.61878329E+01 1.88105120E+00 2.36386368E-02-1.83443295E-05    3
 6.84842963E-09-9.92733674E-13-2.69280190E+04 1.59154793E+01                   4
C2H3OOH    4/18/ 8 THERMC   2H   4O   2    0G   300.000  5000.000 1397.000     1
 1.15749951E+01 8.09909174E-03-2.81808668E-06 4.42697954E-10-2.58998042E-14    2
-8.84852664E+03-3.43859117E+01 1.35644398E+00 3.37002447E-02-2.75988500E-05    3
 1.14222854E-08-1.89488886E-12-5.49996692E+03 1.98354466E+01                   4
C2H3OO                  H   3C   2O   2     G   298.150  2000.000 1000.00      1
 6.04483828E+00 1.45511127E-02-7.50974622E-06 1.83488280E-09-1.66689681E-13    2
 1.01699244E+04-3.71144913E+00 1.09784776E+00 2.95333237E-02-2.27744360E-05    3
 7.20559155E-09-3.07929092E-13 1.13996101E+04 2.13563583E+01                   4
CHCHO                   H   2C   2O   1     G   298.150  2000.000 1000.00      1
 4.92632910E+00 9.71712147E-03-5.54855980E-06 1.53068537E-09-1.64742462E-13    2
 2.89499494E+04 5.27874677E-01 2.33256751E+00 1.62952986E-02-9.72052177E-06    3
 5.15124155E-10 1.03836514E-12 2.96585452E+04 1.39904923E+01                   4
C2H2              G 1/91C  2 H  2    0    0 G   200.000  6000.00  1000.00      1
 4.65878489E+00 4.88396667E-03-1.60828888E-06 2.46974544E-10-1.38605959E-14    2
 2.57594042E+04-3.99838194E+00 8.08679682E-01 2.33615762E-02-3.55172234E-05    3
 2.80152958E-08-8.50075165E-12 2.64289808E+04 1.39396761E+01 2.74459950E+04    4
C2H               T 5/10C  2 H  1    0    0 G   200.000  6000.00  1000.00      1
 3.66270248E+00 3.82492252E-03-1.36632500E-06 2.13455040E-10-1.23216848E-14    2
 6.71683790E+04 3.92205792E+00 2.89867676E+00 1.32988489E-02-2.80733327E-05    3
 2.89484755E-08-1.07502351E-11 6.70616050E+04 6.18547632E+00 6.83210436E+04    4
H2CC              L12/89H   2C   2    0    0G   200.000  6000.000  1000.000    1
 0.42780340E+01 0.47562804E-02-0.16301009E-05 0.25462806E-09-0.14886379E-13    2
 0.48316688E+05 0.64023701E+00 0.32815483E+01 0.69764791E-02-0.23855244E-05    3
-0.12104432E-08 0.98189545E-12 0.48621794E+05 0.59203910E+01 0.49887266E+05    4
C2H5OH     8/12/15      C   2H   6O   1    0G   300.000  5000.000 1402.000     1
 8.14483865E+00 1.28314052E-02-4.29052743E-06 6.55971721E-10-3.76506611E-14    2
-3.24005526E+04-1.86241126E+01 2.15805861E-01 2.95228396E-02-1.68271048E-05    3
 4.49484797E-09-4.02451543E-13-2.94851823E+04 2.45725052E+01                   4
C2H5O      8/12/15      C   2H   5O   1    0G   300.000  5000.000 1467.000     1
 8.19120635E+00 1.10391986E-02-3.75270536E-06 5.80275784E-10-3.35735146E-14    2
-5.66847208E+03-1.90131344E+01 2.90353584E+00 1.77256708E-02-2.69624757E-06    3
-3.45830533E-09 1.25224784E-12-3.28930290E+03 1.13545591E+01                   4
PC2H4OH    8/12/15      C   2H   5O   1    0G   300.000  5000.000 1395.000     1
 8.06750150E+00 1.06143554E-02-3.57999360E-06 5.50363760E-10-3.17051769E-14    2
-6.92747939E+03-1.53833428E+01 2.59479867E+00 2.27100669E-02-1.39473846E-05    3
 4.70095591E-09-6.90044236E-13-4.91486975E+03 1.43240718E+01                   4
SC2H4OH    8/12/15      C   2H   5O   1    0G   300.000  5000.000 1385.000     1
 8.15007136E+00 1.02549305E-02-3.40137764E-06 5.17509965E-10-2.96128942E-14    2
-1.05014386E+04-1.73134615E+01 1.46281093E+00 2.39193995E-02-1.30667185E-05    3
 3.10615465E-09-1.85896007E-13-8.00790323E+03 1.92547092E+01                   4
O2C2H4OH   9/ 1/12 THERMC   2H   5O   3    0G   300.000  5000.000 1506.000     1
 1.27503881E+01 1.11514325E-02-3.83473891E-06 5.98155829E-10-3.48372108E-14    2
-2.52770876E+04-3.54317608E+01 7.04009800E+00 1.59564166E-02 2.21097416E-06    3
-7.05197355E-09 2.08266026E-12-2.24524432E+04-1.75361758E+00                   4
C2H4O2H    9/ 1/12      C   2H   5O   2    0G   300.000  5000.000 1389.000     1
 1.00590614E+01 1.13378955E-02-3.89403387E-06 6.06090687E-10-3.52212353E-14    2
 4.24048653E+02-2.32086536E+01 2.75788364E+00 2.88271987E-02-2.08302264E-05    3
 8.47401397E-09-1.48617610E-12 3.00153893E+03 1.59921711E+01                   4
C2H4O1-2          L 8/88C  2 H  4 O  1    0 G   200.000  6000.00  1000.00      1
 0.54887641E+01 0.12046190E-01-0.43336931E-05 0.70028311E-09-0.41949088E-13    2
-0.91804251E+04-0.70799605E+01 0.37590532E+01-0.94412180E-02 0.80309721E-04    3
-0.10080788E-06 0.40039921E-10-0.75608143E+04 0.78497475E+01-0.63304657E+04    4
C2H3O1-2          A 1/05C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 5.60158035E+00 9.17613962E-03-3.28028902E-06 5.27903888E-10-3.15362241E-14    2
 1.71446252E+04-5.47228512E+00 3.58349017E+00-6.02275805E-03 6.32426867E-05    3
-8.18540707E-08 3.30444505E-11 1.85681353E+04 9.59725926E+00 1.97814471E+04    4
CH3CHO            L 8/88C  2 H  4 O   1   0 G   200.000  6000.00  1000.00      1
 0.54041108E+01 0.11723059E-01-0.42263137E-05 0.68372451E-09-0.40984863E-13    2
-0.22593122E+05-0.34807917E+01 0.47294595E+01-0.31932858E-02 0.47534921E-04    3
-0.57458611E-07 0.21931112E-10-0.21572878E+05 0.41030159E+01-0.19987949E+05    4
CH3CO             IU2/03C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 0.53137165E+01 0.91737793E-02-0.33220386E-05 0.53947456E-09-0.32452368E-13    2
-0.36450414E+04-0.16757558E+01 0.40358705E+01 0.87729487E-03 0.30710010E-04    3
-0.39247565E-07 0.15296869E-10-0.26820738E+04 0.78617682E+01-0.12388039E+04    4
CH2CHO            T03/10C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 6.53928338E+00 7.80238629E-03-2.76413612E-06 4.42098906E-10-2.62954290E-14    2
-1.18858659E+03-8.72091393E+00 2.79502600E+00 1.01099472E-02 1.61750645E-05    3
-3.10303145E-08 1.39436139E-11 1.62944975E+02 1.23646657E+01 1.53380440E+03    4
O2CH2CHO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1393.000     1
 1.11807543E+01 9.14479256E-03-3.15089833E-06 4.91944238E-10-2.86639180E-14    2
-1.55790331E+04-2.87892740E+01-1.29465843E+00 4.44936393E-02-4.26577074E-05    3
 2.07391950E-08-3.96828771E-12-1.18275628E+04 3.60778797E+01                   4
HO2CH2CO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1386.000     1
 1.04146322E+01 1.12680116E-02-5.17494839E-06 1.00333285E-09-6.68165911E-14    2
-1.40955672E+04-2.27894400E+01 2.22681686E+00 3.56781380E-02-3.26401909E-05    3
 1.47651988E-08-2.64794380E-12-1.18735095E+04 1.91581197E+01                   4
C2H3OH     2/ 3/ 9 THERMC   2H   4O   1    0G   300.000  5000.000 1410.000     1
 8.32598158E+00 8.03387281E-03-2.63928405E-06 3.98410726E-10-2.26551155E-14    2
-1.83221436E+04-2.02080305E+01-1.27972260E-01 3.38506073E-02-3.30644935E-05    3
 1.64858739E-08-3.19935455E-12-1.59914544E+04 2.30438601E+01                   4
C2H2OH                  H   3C   2O   1    0G   300.000  5000.000 1401.000     1
 8.20268447E+00 5.92989165E-03-1.99194448E-06 3.05794341E-10-1.76114732E-14    2
 1.24881328E+04-1.89670436E+01 6.41642616E-01 2.61903633E-02-2.30385370E-05    3
 1.02804704E-08-1.81971416E-12 1.48276951E+04 2.06750999E+01                   4
CH2CO                   H   2C   2O   1    0G    300.00   5000.00 1000.00      1
 5.35869367E+00 6.95641586E-03-2.64802637E-06 4.65067592E-10-3.08641820E-14    2
-7.90294013E+03-3.98525731E+00 1.81422511E+00 1.99008590E-02-2.21416008E-05    3
 1.45028521E-08-3.98877068E-12-7.05394926E+03 1.36079359E+01                   4
HCCO              T 4/09H  1 C  2 O  1    0 G   200.000  6000.00  1000.00      1
 5.91479333E+00 3.71408730E-03-1.30137010E-06 2.06473345E-10-1.21476759E-14    2
 1.93596301E+04-5.50567269E+00 1.87607969E+00 2.21205418E-02-3.58869325E-05    3
 3.05402541E-08-1.01281069E-11 2.01633840E+04 1.36968290E+01 2.14444387E+04    4
HCCOH             T12/09C  2 H  2 O  1    0 G   200.000  6000.00  1000.00      1
 6.37509678E+00 5.49429011E-03-1.88136576E-06 2.93803536E-10-1.71771901E-14    2
 8.93277676E+03-8.24498007E+00 2.05541154E+00 2.52003372E-02-3.80821654E-05    3
 3.09890632E-08-9.89799902E-12 9.76872113E+03 1.22271534E+01 1.12217316E+04    4
CH3CO3H    6/26/95 THERMC   2H   4O   3    0G   300.000  5000.000 1391.000     1
 1.25060485E+01 9.47789695E-03-3.30402246E-06 5.19630793E-10-3.04233568E-14    2
-4.59856703E+04-3.79195947E+01 2.24135876E+00 3.37963514E-02-2.53887482E-05    3
 9.67583587E-09-1.49266157E-12-4.24677831E+04 1.70668133E+01                   4
CH3CO3     4/ 3/ 0 THERMC   2H   3O   3    0G   300.000  5000.000 1391.000     1
 1.12522498E+01 8.33652672E-03-2.89014530E-06 4.52781734E-10-2.64354456E-14    2
-2.60238584E+04-2.96370457E+01 3.60373432E+00 2.70080341E-02-2.08293438E-05    3
 8.50541104E-09-1.43846110E-12-2.34205171E+04 1.12014914E+01                   4
CH3CO2     2/14/95 THERMC   2H   3O   2    0G   300.000  5000.000 1395.000     1
 8.54059736E+00 8.32951214E-03-2.84722010E-06 4.41927196E-10-2.56373394E-14    2
-2.97290678E+04-2.03883545E+01 1.37440768E+00 2.49115604E-02-1.74308894E-05    3
 6.24799508E-09-9.09516835E-13-2.72330150E+04 1.81405454E+01                   4
CH3OCH3    2/11/14 THERMC   2H   6O   1    0G   300.000  5000.000 1999.000     1
 6.03232751E+00 1.56155270E-02-5.50761030E-06 8.75666140E-10-5.17180562E-14    2
-2.52690354E+04-8.25885183E+00 2.05597390E+00 2.07019456E-02-5.00382376E-06    3
-1.62279885E-09 6.84330155E-13-2.35494445E+04 1.45029944E+01                   4
CH3OCH2    2/11/14 THERMC   2H   5O   1    0G   300.000  5000.000 1395.000     1
 6.62621974E+00 1.22219496E-02-4.12416696E-06 6.34127512E-10-3.65317390E-14    2
-3.33965890E+03-8.95305753E+00 1.58874948E+00 2.24414123E-02-1.19434933E-05    3
 3.37160213E-09-4.15077249E-13-1.37208255E+03 1.87548958E+01                   4
CH3OCH2O2H 2/12/14 THERMC   2H   6O   3    0G   300.000  5000.000 1404.000     1
 1.28159161E+01 1.34818095E-02-4.50397729E-06 6.88229286E-10-3.94883680E-14    2
-4.06745921E+04-3.78047802E+01 1.05786981E+00 4.36787095E-02-3.46383899E-05    3
 1.44808830E-08-2.46100643E-12-3.68851076E+04 2.43391936E+01                   4
CH3OCH2O2  2/12/14 THERMC   2H   5O   3    0G   300.000  5000.000 1441.000     1
 1.19179361E+01 1.19412867E-02-3.93526185E-06 5.95756132E-10-3.39597705E-14    2
-2.34231833E+04-3.20096863E+01 3.39930541E+00 3.09460407E-02-1.92548181E-05    3
 5.76033887E-09-6.16081571E-13-2.04433218E+04 1.39429608E+01                   4
CH2OCH2O2H 2/12/14 THERMC   2H   5O   3    0G   300.000  5000.000 1418.000     1
 1.23892901E+01 1.11758961E-02-3.59249095E-06 5.34196366E-10-3.00536541E-14    2
-1.80551598E+04-3.29576862E+01 1.62245477E-01 4.76101093E-02-4.52046954E-05    3
 2.18379311E-08-4.11295947E-12-1.46498100E+04 2.98253164E+01                   4
O2CH2OCH2O2H 2/12/14 ERMC   2H   5O   5    0G   300.000  5000.000 1433.000     1
 1.77378326E+01 1.13589899E-02-3.67382539E-06 5.49255712E-10-3.10405899E-14    2
-3.82903058E+04-5.66609932E+01 2.39977678E+00 5.39881943E-02-4.87969524E-05    3
 2.19792134E-08-3.86106979E-12-3.37824638E+04 2.30683371E+01                   4
HO2CH2OCHO 2/12/14 THERMC   2H   4O   4    0G   300.000  5000.000 1386.000     1
 1.57136128E+01 9.64430166E-03-3.44136025E-06 5.49722196E-10-3.25360322E-14    2
-6.29409094E+04-5.29505242E+01 1.21909586E+00 4.28858235E-02-3.17634222E-05    3
 1.11542676E-08-1.49753153E-12-5.79287926E+04 2.49759193E+01                   4
OCH2OCHO   5/29/14 THERMC   2H   3O   3    0G   300.000  5000.000 1523.000     1
 1.24013200E+01 7.83738243E-03-2.82992688E-06 4.55558739E-10-2.71061389E-14    2
-4.68453470E+04-3.78084549E+01 1.89539692E+00 2.74118545E-02-1.36476090E-05    3
 1.26325603E-09 5.17970476E-13-4.27879440E+04 2.02333278E+01                   4
HOCH2OCO   5/29/14 THERMC   2H   3O   3    0G   300.000  5000.000 1443.000     1
 1.11498410E+01 9.34736520E-03-3.35541548E-06 5.38037115E-10-3.19260183E-14    2
-4.75012119E+04-2.95983867E+01 5.95255071E+00 8.42196282E-03 1.36741678E-05    3
-1.46786275E-08 3.84143533E-12-4.44470269E+04 2.85657217E+00                   4
CH3OCH2O   5/15/14 THERMC   2H   5O   2    0G   300.000  5000.000 1523.000     1
 9.81288609E+00 1.21313106E-02-4.30285768E-06 6.84443177E-10-4.03862658E-14    2
-2.50760742E+04-2.51866352E+01 5.63414373E+00 8.92830283E-03 1.37225633E-05    3
-1.40497059E-08 3.54625624E-12-2.22825214E+04 1.93588846E+00                   4
CH3OCHO           T 6/08C  2 H  4 O  2    0 G   200.000  6000.00  1000.00      1
 6.33360880E+00 1.34851485E-02-4.84305805E-06 7.81719241E-10-4.67917447E-14    2
-4.68316521E+04-6.91542601E+00 5.96757028E+00-9.38085425E-03 7.07648417E-05    3
-8.29932227E-08 3.13522917E-11-4.55713267E+04 7.50341113E-01-4.37330508E+04    4
CH3OCO     5/ 8/ 3 THERMC   2H   3O   2    0G   300.000  5000.000 1601.000     1
 9.73659803E+00 7.42432713E-03-2.65641779E-06 4.25031143E-10-2.51824924E-14    2
-2.36015721E+04-2.36353471E+01 4.16215406E+00 1.38037511E-02-3.08486109E-07    3
-4.56430814E-09 1.46909632E-12-2.10130301E+04 8.64301044E+00                   4
CH2OCHO    4/15/ 8 THERMC   2H   3O   2    0G   300.000  5000.000 1442.000     1
 1.00960096E+01 7.19887066E-03-2.59813465E-06 4.18110812E-10-2.48723387E-14    2
-2.36389018E+04-2.71144175E+01 2.31031671E+00 1.80474065E-02-2.71519637E-06    3
-4.60918579E-09 1.70037078E-12-2.02910878E+04 1.71549722E+01                   4
C3H8       8/12/15      C   3H   8    0    0G   300.000  5000.000 1390.000     1
 9.15541310E+00 1.72574139E-02-5.85614868E-06 9.04190155E-10-5.22523772E-14    2
-1.75762439E+04-2.77418510E+01 2.40878470E-01 3.39548599E-02-1.60930874E-05    3
 2.83480628E-09 2.78195172E-14-1.40362853E+04 2.16500800E+01                   4
IC3H7      8/12/15      C   3H   7    0    0G   298.000  6000.0    1000.0      1
 6.70775549E+00 1.74048076E-02-6.07615926E-06 9.60084351E-10-5.65656490E-14    2
 7.55377821E+03-1.03686516E+01-8.97467137E-01 4.15744022E-02-4.94778349E-05    3
 4.56493655E-08-1.79085437E-11 9.93950407E+03 2.92641758E+01                   4
NC3H7      8/12/15      C   3H   7    0    0G   298.0    6000.0    1000.0      1
 7.48614243E+00 1.65769478E-02-5.74876481E-06 9.04103694E-10-5.30867231E-14    2
 8.93710008E+03-1.42595379E+01-2.20120865E+00 5.29641653E-02-7.23640506E-05    3
 6.36996940E-08-2.29332581E-11 1.15130744E+04 3.43669174E+01                   4
NC3H7O2H   8/12/15      C   3H   8O   2    0G   300.000  5000.000 1392.000     1
 1.42246236E+01 1.74340964E-02-5.97063522E-06 9.27753851E-10-5.38585168E-14    2
-2.88159737E+04-4.74357865E+01 1.35815897E+00 4.56683952E-02-2.91646368E-05    3
 9.41701313E-09-1.22337394E-12-2.41528416E+04 2.23322825E+01                   4
NC3H7O2    8/12/15      C   3H   7O   2    0G   300.000  5000.000 1390.000     1
 1.32753283E+01 1.61303126E-02-5.52348308E-06 8.58197168E-10-4.98172586E-14    2
-1.16032968E+04-4.15091215E+01 2.13311681E+00 3.96692045E-02-2.37570127E-05    3
 6.96020417E-09-7.82576856E-13-7.46687112E+03 1.92444565E+01                   4
IC3H7O2H   8/12/15      C   3H   8O   2    0G   300.000  5000.000 1405.000     1
 1.44896107E+01 1.68268026E-02-5.67601391E-06 8.72850837E-10-5.02993991E-14    2
-3.06478491E+04-5.01352281E+01 1.77384705E+00 4.75813498E-02-3.43745304E-05    3
 1.31405381E-08-2.06922904E-12-2.63458844E+04 1.77669753E+01                   4
IC3H7O2    8/12/15      C   3H   7O   2    0G   300.000  5000.000 1407.000     1
 1.35268120E+01 1.54306581E-02-5.17464218E-06 7.92548669E-10-4.55415379E-14    2
-1.33946348E+04-4.40461451E+01 2.58517502E+00 4.16107259E-02-2.92193877E-05    3
 1.08614807E-08-1.66312005E-12-9.67013161E+03 1.44731300E+01                   4
NC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1386.000     1
 1.15279177E+01 1.53775991E-02-5.23946272E-06 8.11382512E-10-4.69927603E-14    2
-9.85099867E+03-3.54233008E+01 2.57486880E+00 3.07100600E-02-1.20048836E-05    3
 3.40807108E-12 7.25275283E-13-6.20913350E+03 1.45966401E+01                   4
IC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1527.000     1
 1.19648494E+01 1.42943974E-02-4.71413211E-06 7.14027066E-10-4.07161162E-14    2
-1.17519389E+04-3.88860959E+01 2.36108410E+00 3.45650027E-02-1.94579631E-05    3
 4.71536901E-09-2.64704937E-13-8.28791395E+03 1.33112436E+01                   4
C3H6OOH1-2 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1387.000     1
 1.38088686E+01 1.43845650E-02-4.74440961E-06 7.19308280E-10-4.10654123E-14    2
-5.14352831E+03-4.20210765E+01 2.83631132E+00 3.88229894E-02-2.47944364E-05    3
 7.85644898E-09-9.58634300E-13-1.26002528E+03 1.72549973E+01                   4
C3H6OOH1-3 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1401.000     1
 1.39130757E+01 1.40218463E-02-4.55921149E-06 6.84182417E-10-3.87696213E-14    2
-3.65650518E+03-4.21532559E+01 1.74271107E+00 4.53733504E-02-3.57580373E-05    3
 1.48540053E-08-2.49981756E-12 2.32580844E+02 2.20973041E+01                   4
C3H6OOH2-1 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1393.000     1
 1.36645362E+01 1.54329764E-02-5.29285952E-06 8.23001262E-10-4.77931121E-14    2
-5.58295862E+03-4.28758364E+01 2.38465746E+00 4.42928555E-02-3.50977087E-05    3
 1.53695144E-08-2.81167824E-12-1.80979612E+03 1.69923285E+01                   4
C3H6OOH1-2O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1404.000     1
 1.91044980E+01 1.44076100E-02-4.72127814E-06 7.12631642E-10-4.05578490E-14    2
-2.50270510E+04-6.63747978E+01 3.99085043E+00 5.31865338E-02-4.28597948E-05    3
 1.77187019E-08-2.92768695E-12-2.02143526E+04 1.34150719E+01                   4
C3H6OOH1-3O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1416.000     1
 1.81661664E+01 1.47644887E-02-4.74842743E-06 7.06972467E-10-3.98305587E-14    2
-2.26256376E+04-5.93719393E+01 5.56933350E+00 4.68523421E-02-3.58917784E-05    3
 1.43314525E-08-2.29776083E-12-1.86065694E+04 7.18655005E+00                   4
C3H6OOH2-1O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1404.000     1
 1.91044980E+01 1.44076100E-02-4.72127814E-06 7.12631642E-10-4.05578490E-14    2
-2.50270510E+04-6.63747978E+01 3.99085043E+00 5.31865338E-02-4.28597948E-05    3
 1.77187019E-08-2.92768695E-12-2.02143526E+04 1.34150719E+01                   4
C3KET12   10/17/12      C   3H   6O   3    0G   300.000  5000.000 1385.000     1
 1.70187760E+01 1.32097361E-02-4.67054741E-06 7.41411770E-10-4.36869787E-14    2
-4.23572589E+04-5.92615939E+01 1.03882879E+00 5.34180080E-02-4.47684141E-05    3
 1.94651680E-08-3.45055244E-12-3.70308881E+04 2.56511209E+01                   4
C3KET13   10/17/12      C   3H   6O   3    0G   300.000  5000.000 1508.000     1
 1.73612692E+01 1.32330813E-02-4.75332110E-06 7.62529227E-10-4.52613717E-14    2
-4.06248060E+04-6.17768199E+01 4.74956819E+00 3.14080991E-02-6.83838427E-06    3
-5.67123901E-09 2.27686972E-12-3.51924570E+04 9.83753744E+00                   4
C3H51-2,3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1386.000     1
 2.12378169E+01 1.39519596E-02-4.94539222E-06 7.86381389E-10-4.63925564E-14    2
-1.92864584E+04-7.69636561E+01 2.55619708E+00 6.13504487E-02-5.23205391E-05    3
 2.28208029E-08-4.02231508E-12-1.31353414E+04 2.21043799E+01                   4
C3H52-1,3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1379.000     1
 2.02817964E+01 1.48155431E-02-5.25503386E-06 8.35963453E-10-4.93308915E-14    2
-1.80085066E+04-7.22688262E+01 4.12253742E+00 5.19553611E-02-3.83733727E-05    3
 1.45851637E-08-2.29820536E-12-1.22759164E+04 1.48367359E+01                   4
C3H5O1-2OOH-3 10/13 THERC   3H   6O   3    0G   300.000  5000.000 1432.000     1
 1.57042382E+01 1.30255692E-02-4.23544254E-06 6.35555595E-10-3.60110207E-14    2
-2.77269333E+04-5.51895464E+01-3.25001215E+00 6.65787151E-02-6.18859778E-05    3
 2.84638649E-08-5.08511634E-12-2.22371240E+04 4.30381280E+01                   4
C3H5O1-3OOH-2 10/13 THERC   3H   6O   3    0G   300.000  5000.000 1434.000     1
 1.44493479E+01 1.36372560E-02-4.25836513E-06 6.20006211E-10-3.43451580E-14    2
-2.77372360E+04-5.06099103E+01-4.43959178E+00 7.16532928E-02-7.15032351E-05    3
 3.51737842E-08-6.63682938E-12-2.27250412E+04 4.56394038E+01                   4
C3H6O1-2          A01/05C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 8.01491079E+00 1.73919953E-02-6.26027968E-06 1.01188256E-09-6.06239111E-14    2
-1.51980838E+04-1.88279964E+01 3.42806676E+00 6.25176642E-03 6.13196311E-05    3
-8.60387185E-08 3.51371393E-11-1.28446646E+04 1.04244994E+01-1.11564001E+04    4
C3H6O1-3          A11/04C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 6.80716906E+00 1.88824545E-02-6.79082475E-06 1.09713919E-09-6.57154952E-14    2
-1.36547629E+04-1.35382154E+01 5.15283752E+00-1.86401716E-02 1.29980652E-04    3
-1.58629974E-07 6.20668783E-11-1.13243512E+04 4.73561224E+00-9.75233898E+03    4
C3H6       8/12/15      C   3H   6    0    0G   298.000  6000.000 1000.000     1
 6.59032304E+00 1.52592866E-02-5.30369441E-06 8.35510888E-10-4.91215549E-14    2
-2.47481113E+02-1.15748238E+01-1.54606737E+00 4.36553128E-02-5.61392417E-05    3
 4.98421927E-08-1.84798923E-11 2.07056233E+03 2.99232495E+01                   4
C3H5-A     8/12/15      C   3H   5    0    0G   298.000  6000.000 1000.000     1
 7.37604097E+00 1.23449782E-02-4.26463882E-06 6.69045835E-10-3.92202554E-14    2
 1.77332960E+04-1.61758204E+01-3.32899442E+00 5.38423469E-02-7.65500752E-05    3
 6.35512285E-08-2.14283003E-11 2.03420628E+04 3.68038362E+01                   4
C3H5-S     8/12/15      C   3H   5    0    0G   300.000  5000.000 1390.000     1
 7.95954498E+00 1.11163183E-02-3.75197834E-06 5.77246260E-10-3.32768957E-14    2
 2.80567891E+04-1.79800372E+01 1.61793372E+00 2.44803904E-02-1.41856503E-05    3
 4.16402233E-09-4.90904795E-13 3.04291037E+04 1.66341443E+01                   4
C3H5-T     8/12/15      C   3H   5    0    0G   300.000  5000.000 1376.000     1
 7.69949212E+00 1.17803985E-02-4.07791749E-06 6.38119222E-10-3.72229675E-14    2
 2.61747145E+04-1.68305890E+01 2.29256998E+00 1.98527646E-02-6.42635654E-06    3
-5.90016395E-10 5.05491095E-13 2.85773377E+04 1.39407124E+01                   4
CC3H6                   C   3H   6O   0    0G   200.000  6000.000 1000.        1
 6.21663437E+00 1.65393591E-02-5.90075838E-06 9.48095199E-10-5.65661522E-14    2
 2.95937491E+03-1.36041009E+01 2.83278674E+00-5.21028618E-03 9.29583210E-05    3
-1.22753194E-07 4.99191366E-11 5.19520048E+03 1.08306333E+01 6.41047999E+03    4
C3H5O             KPS12 C   3H   5O   1    0G   300.000  5000.000 1402.000     1
 1.02638186E+01 1.17609932E-02-3.89837957E-06 5.92650815E-10-3.38867417E-14    2
 7.25938472E+03-2.75108651E+01 8.24068673E-01 3.46749909E-02-2.51786795E-05    3
 9.56781953E-09-1.48085302E-12 1.04203725E+04 2.28283070E+01                   4
CH2CHOCH2  8/ 8/15      C   3H   5O   1    0G   300.000  5000.000 1384.000     1
 1.20076931E+01 1.05055204E-02-3.69920541E-06 5.85629983E-10-3.44431587E-14    2
 6.97311613E+03-3.75189859E+01 1.15350351E+00 3.51253596E-02-2.50071619E-05    3
 9.00715632E-09-1.32376643E-12 1.08300872E+04 2.10606652E+01                   4
CH3CHCHO                C   3H   5O   1    0G   300.000  5000.000 1424.000     1
 1.06781476E+01 1.12805711E-02-3.89010759E-06 6.07617268E-10-3.54120848E-14    2
-7.73234209E+03-3.24971238E+01 1.47166733E+00 2.69251618E-02-1.00248013E-05    3
-1.13421435E-09 1.03416658E-12-4.04142023E+03 1.88722472E+01                   4
AC4H7OOH   6/17/13 THERMC   4H   8O   2    0G   300.000  5000.000 1395.000     1
 1.47661443E+01 2.12235231E-02-7.09403390E-06 1.08423759E-09-6.22145708E-14    2
-1.35617411E+04-4.77449138E+01 1.33470633E+00 5.27831440E-02-3.58861360E-05    3
 1.32495013E-08-2.06619289E-12-8.87891782E+03 2.43857336E+01                   4
C3H6OH1-2  9/ 1/12      C   3H   7O   1    0G   300.000  5000.000 1395.000     1
 1.00338281E+01 1.60227373E-02-5.41658448E-06 8.34191172E-10-4.81215988E-14    2
-1.27912397E+04-2.39034395E+01 5.05207596E-01 3.63869988E-02-2.15530901E-05    3
 6.45584786E-09-7.71267046E-13-9.26980840E+03 2.79804349E+01                   4
CH3CHCO   03/03/95 THERMC   3H   4O   1    0G   300.000  5000.000 1400.00      1
 1.00219123E+01 9.56966300E-03-3.26221644E-06 5.05231706E-10-2.92593257E-14    2
-1.42482738E+04-2.77829973E+01 1.48380119E+00 3.22203013E-02-2.70250033E-05    3
 1.20499164E-08-2.18365931E-12-1.15276540E+04 1.71552068E+01                   4
AC3H5OOH    GOLDSMITH   C   3H   6O   2    0G   298.0    6000.0   1000.000     1
 1.20838649E+01 1.47946591E-02-5.13212591E-06 8.07504999E-10-4.74394983E-14    2
-1.02184463E+04-3.36434791E+01 3.18124993E+00 4.35233041E-02-5.16277353E-05    3
 4.32011427E-08-1.57714983E-11-7.63521503E+03 1.21725683E+01                   4
C3H6OH2-1  8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000     1
 1.12222277E+01 1.36444398E-02-4.51406709E-06 7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01 1.09670360E+00 3.80727565E-02-2.75022497E-05    3
 1.07477493E-08-1.74895773E-12-1.40764487E+04 2.22475799E+01                   4
HOC3H6O2   9/ 1/12      C   3H   7O   3    0G   300.000  5000.000 1407.000     1
 1.56948113E+01 1.57703692E-02-5.30501726E-06 8.14307835E-10-4.68666193E-14    2
-3.24540840E+04-5.06084117E+01 2.84960487E+00 4.77244552E-02-3.60392974E-05    3
 1.43479922E-08-2.33507634E-12-2.82106103E+04 1.76478537E+01                   4
SC3H5OH    2/ 3/ 9      C   3H   6O   1    0G   300.000  5000.000 1404.000     1
 1.11222064E+01 1.27745410E-02-4.25315532E-06 6.48216484E-10-3.71190850E-14    2
-2.36690795E+04-3.41335182E+01-3.53977226E-02 4.34969453E-02-3.74479918E-05    3
 1.70906074E-08-3.13775054E-12-2.02502608E+04 2.41528201E+01                   4
IC3H5OH    8/ 1/95 THERMC   3H   6O   1    0G   300.000  5000.000 1374.00      1
 1.07381025E+01 1.31698194E-02-4.41529622E-06 6.77009837E-10-3.89608901E-14    2
-2.47298321E+04-3.13634050E+01 1.58376391E+00 3.16215366E-02-1.73664942E-05    3
 4.18927663E-09-2.79899620E-13-2.12643496E+04 1.88313766E+01                   4
C3H5OH            T06/10C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 8.72477114E+00 1.63942712E-02-5.90852993E-06 9.53262253E-10-5.70318010E-14    2
-1.90496618E+04-1.97198674E+01 3.15011905E+00 1.28538274E-02 4.28438434E-05    3
-6.67818707E-08 2.80408237E-11-1.66413668E+04 1.35066359E+01-1.48710589E+04    4
CH2CCH2OH  9/ 8/95 THERMC   3H   5O   1    0G   300.000  5000.000 1372.00      1
 9.70702027E+00 1.13972660E-02-3.77993962E-06 5.75209277E-10-3.29229125E-14    2
 9.13212884E+03-2.25012933E+01 2.88422544E+00 2.42428071E-02-1.14152268E-05    3
 1.71775334E-09 1.42177454E-13 1.17935615E+04 1.52102335E+01                   4
C3H4-P            T 2/90H  4 C  3    0    0 G   200.000  6000.00  1000.00      1
 0.60252400E+01 0.11336542E-01-0.40223391E-05 0.64376063E-09-0.38299635E-13    2
 0.19620942E+05-0.86043785E+01 0.26803869E+01 0.15799651E-01 0.25070596E-05    3
-0.13657623E-07 0.66154285E-11 0.20802374E+05 0.98769351E+01 0.22302059E+05    4
C3H4-A            L 8/89C  3 H  4    0    0 G   200.000  6000.00  1000.00      1
 0.63168722E+01 0.11133728E-01-0.39629378E-05 0.63564238E-09-0.37875540E-13    2
 0.20117495E+05-0.10995766E+02 0.26130445E+01 0.12122575E-01 0.18539880E-04    3
-0.34525149E-07 0.15335079E-10 0.21541567E+05 0.10226139E+02 0.22962267E+05    4
C3H3              T 7/11C  3 H  3    0    0 G   200.000  6000.00  1000.000     1
 7.14221719E+00 7.61902211E-03-2.67460030E-06 4.24914904E-10-2.51475443E-14    2
 3.95709594E+04-1.25848690E+01 1.35110873E+00 3.27411291E-02-4.73827407E-05    3
 3.76310220E-08-1.18541128E-11 4.07679941E+04 1.52058598E+01 4.22762135E+04    4
CC3H4             T12/81C   3H   4    0    0G   300.000  5000.00  1000.00      1
 0.66999931E+01 0.10357372E-01-0.34551167E-05 0.50652949E-09-0.26682276E-13    2
 0.30199051E+05-0.13378770E+02-0.24621047E-01 0.23197215E-01-0.18474357E-05    3
-0.15927593E-07 0.86846155E-11 0.32334137E+05 0.22729762E+02 0.33327280E+05    4
C3H2              T12/00C  3 H  2    0    0 G   200.000  6000.00  1000.00      1
 6.67324762E+00 5.57728845E-03-1.99180164E-06 3.20289156E-10-1.91216272E-14    2
 7.57571184E+04-9.72894405E+00 2.43417332E+00 1.73013063E-02-1.18294047E-05    3
 1.02756396E-09 1.62626314E-12 7.69074892E+04 1.21012230E+01 7.83005132E+04    4
H2CCC(S)               0C   3H   2    0    0G   200.000  5000.000 1500.00      1
 0.64888762E+01 0.53112789E-02-0.17809490E-05 0.27252642E-09-0.15619590E-13    2
 0.63661864E+05-0.10064283E+02 0.37229726E+01 0.92589854E-02-0.23006191E-05    3
-0.10200808E-08 0.45374357E-12 0.64877289E+05 0.56865936E+01                   4
C3H2(S)                0C   3H   2    0    0G   200.000  5000.000  900.00      1
 0.77642570E+01 0.47112774E-02-0.16170637E-05 0.25472406E-09-0.15038572E-13    2
 0.66849672E+05-0.15098549E+02 0.52976482E+01 0.16987466E-01-0.24266517E-04    3
 0.18653681E-07-0.55763001E-11 0.67240466E+05-0.37540041E+01                   4
C3H2C                  0C   3H   2    0    0G   200.000  5000.000 1500.00      1
 0.65632680E+01 0.52363256E-02-0.17544830E-05 0.26866106E-09-0.15428509E-13    2
 0.56514618E+05-0.12000607E+02 0.11295888E+01 0.17287401E-01-0.11366823E-04    3
 0.34569296E-08-0.36615951E-12 0.58419080E+05 0.17331448E+02                   4
PC3H4OH-2  4/ 2/13 THERMC   3H   5O   1    0G   300.000  5000.000 1403.000     1
 1.07164095E+01 1.06066461E-02-3.51374060E-06 5.33713932E-10-3.04901511E-14    2
 4.98486803E+03-2.98329329E+01 1.42757363E+00 3.64825569E-02-3.18007132E-05    3
 1.46914605E-08-2.72331227E-12 7.80342663E+03 1.85890339E+01                   4
SC3H4OH    3/28/13      C   3H   5O   1    0G   300.000  5000.000 1407.000     1
 1.20968484E+01 9.43976596E-03-3.10773897E-06 4.69609188E-10-2.67165710E-14    2
-3.85854894E+02-3.76795997E+01 1.72870561E+00 4.41015870E-02-4.72013860E-05    3
 2.52073596E-08-5.13375710E-12 2.22720503E+03 1.43928257E+01                   4
C3H3O      2/17/14 CZHOUH   3C   3O   1     G   298.150  2000.000 1000.00      1
 4.19355696E+00 1.95625103E-02-1.22336450E-05 3.90615061E-09-5.08539231E-13    2
 3.14931737E+04 5.03216224E+00 8.75023836E-01 3.51184068E-02-3.89901356E-05    3
 2.40255750E-08-6.10883631E-12 3.20427921E+04 2.04717253E+01                   4
C3H3O2H    1/31/13      C   3H   4O   2    0G   300.000  5000.000 1385.000     1
 1.38152174E+01 8.62174763E-03-3.06710006E-06 4.88874247E-10-2.88888385E-14    2
 6.29182941E+03-4.39151257E+01 1.09787313E+00 4.22717882E-02-3.83969355E-05    3
 1.77405069E-08-3.27674312E-12 1.03592314E+04 2.30651783E+01                   4
C2HCHO     1/31/13      C   3H   2O   1    0G   300.000  5000.000 2012.000     1
 7.99952054E+00 7.07825497E-03-2.63086819E-06 4.33073185E-10-2.62003284E-14    2
 8.71863156E+03-1.57226237E+01 4.20776611E+00 1.34382727E-02-5.15442099E-06    3
-2.24570818E-11 2.74111284E-13 1.02117375E+04 5.43871873E+00                   4
C2H5CHO    8/12/15      C   3H   6O   1    0G   300.000  5000.000 1449.000     1
 1.06224453E+01 1.35569132E-02-4.60754771E-06 7.12755462E-10-4.12631683E-14    2
-2.78692266E+04-3.16628752E+01 2.18895588E+00 2.58289987E-02-6.04170058E-06    3
-3.70702654E-09 1.57131095E-12-2.42671146E+04 1.61496330E+01                   4
C2H5CO            A10/04C  3 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 6.52325448E+00 1.54211952E-02-5.50898157E-06 8.85889862E-10-5.28846399E-14    2
-7.19631634E+03-5.19862218E+00 6.25722402E+00-9.17612184E-03 7.61190493E-05    3
-9.05514997E-08 3.46198215E-11-5.91616484E+03 2.23330599E+00-3.94851891E+03    4
CH2CH2CHO               C   3H   5O   1    0G   300.000  5000.000 1437.000     1
 1.00673122E+01 1.14971005E-02-3.90137798E-06 6.03029101E-10-3.48958224E-14    2
-2.75080876E+03-2.58818404E+01 2.55799036E+00 2.23391941E-02-4.89741478E-06    3
-3.58874384E-09 1.47175030E-12 4.53127696E+02 1.67016285E+01                   4
C2H3CHO           KPS12 C   3H   4O   1    0G   300.000  5000.000 1398.000     1
 9.99155394E+00 9.82348001E-03-3.31203088E-06 5.09524422E-10-2.93821890E-14    2
-1.25303509E+04-2.85168883E+01 7.33844455E-01 3.17482671E-02-2.29599468E-05    3
 8.42104232E-09-1.23613478E-12-9.38473548E+03 2.10308851E+01                   4
C2H3CO            KPS12 C   3H   3O   1    0G   300.000  5000.000 1395.000     1
 8.86032735E+00 8.48985205E-03-2.90350080E-06 4.50763986E-10-2.61524281E-14    2
 7.73489171E+03-2.06978792E+01 1.65335195E+00 2.57402596E-02-1.89009911E-05    3
 7.29174972E-09-1.16083226E-12 1.02020654E+04 1.78705872E+01                   4
CH3COCH3   8/12/15      C   3H   6O   1    0G   300.000  5000.000 1394.000     1
 8.87619308E+00 1.45700263E-02-4.84823280E-06 7.38614777E-10-4.22831194E-14    2
-3.06046242E+04-2.12730484E+01 2.20008426E+00 2.74019559E-02-1.31342003E-05    3
 2.57150371E-09-6.21509091E-14-2.79933966E+04 1.55883508E+01                   4
CH3COCH2   2/14/13 THERMC   3H   5O   1    0G   300.000  5000.000 1387.000     1
 1.09524298E+01 1.11458668E-02-3.86262877E-06 6.05088857E-10-3.53293362E-14    2
-9.60833727E+03-3.15622776E+01 1.13381826E+00 3.25095045E-02-2.10424651E-05    3
 6.64421151E-09-8.12618901E-13-6.04868361E+03 2.17158655E+01                   4
CH3COCH2O2 2/14/13 THERMC   3H   5O   3    0G   300.000  5000.000 1397.000     1
 1.65756401E+01 1.06465489E-02-3.61368681E-06 5.59053564E-10-3.23832271E-14    2
-2.42541401E+04-5.45304899E+01 1.19378141E+00 4.98027161E-02-4.17999508E-05    3
 1.74527607E-08-2.88198761E-12-1.93244224E+04 2.67877493E+01                   4
CH3COCH2O  2/ 8/13 THERMC   3H   5O   2    0G   300.000  5000.000 2002.000     1
 9.84061707E+00 1.59181106E-02-5.85164644E-06 9.56160073E-10-5.75477263E-14    2
-2.11214823E+04-2.12330791E+01 5.85960137E+00 1.78954926E-02 7.41506398E-07    3
-5.40032753E-09 1.47393197E-12-1.90714739E+04 2.70987883E+00                   4
C3KET21    2/14/13 THERMC   3H   6O   3    0G   300.000  5000.000 1394.000     1
 1.75768076E+01 1.20311704E-02-4.11633942E-06 6.40149366E-10-3.72127562E-14    2
-4.15502347E+04-6.09097100E+01-8.74352903E-01 6.12501498E-02-5.51474542E-05    3
 2.48491014E-08-4.42613472E-12-3.58060819E+04 3.59306224E+01                   4
C4H10      8/12/15      C   4H  10    0    0G   300.000  5000.000 1392.000     1
 1.24923813E+01 2.15951935E-02-7.34277611E-06 1.13529859E-09-6.56730149E-14    2
-2.17598985E+04-4.41546866E+01-9.20862487E-02 4.69703816E-02-2.54761945E-05    3
 6.35894738E-09-5.16005946E-13-1.69556758E+04 2.49101571E+01                   4
PC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1393.000     1
 1.18547949E+01 1.96962095E-02-6.71054229E-06 1.03891144E-09-6.01513573E-14    2
 3.38182243E+03-3.72343446E+01 4.09644702E-01 4.29511341E-02-2.36582809E-05    3
 6.15744917E-09-5.64300671E-13 7.74319150E+03 2.55312526E+01                   4
SC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1682.000     1
 9.25139144E+00 2.24301385E-02-7.82648592E-06 1.23559460E-09-7.26249864E-14    2
 3.11148804E+03-2.16080436E+01 9.42662332E-01 3.77414530E-02-1.58911963E-05    3
 1.75489317E-09 2.89725750E-13 6.20542636E+03 2.42126605E+01                   4
PC4H9O                  C   4H   9O   1    0G   300.000  5000.000 1396.000     1
 1.53371588E+01 1.92789649E-02-6.56856538E-06 1.01724003E-09-5.89183466E-14    2
-1.41958782E+04-5.45071855E+01 1.84659093E+00 4.61054365E-02-2.44856516E-05    3
 5.11293268E-09-1.07538298E-13-9.09206746E+03 1.95237441E+01                   4
SC4H9O                  C   4H   9O   1    0G   300.000  5000.000 1411.000     1
 1.52130012E+01 1.90029969E-02-6.39004701E-06 9.80774402E-10-5.64493733E-14    2
-1.59888805E+04-5.43195369E+01 2.01772535E+00 4.70083969E-02-2.74726645E-05    3
 7.36290028E-09-6.30414237E-13-1.11892176E+04 1.74371746E+01                   4
PC4H9O2    8/12/15      C   4H   9O   2    0G   300.000  5000.000 1391.000     1
 1.66120049E+01 2.04752336E-02-7.01415262E-06 1.09010510E-09-6.32913959E-14    2
-1.57901735E+04-5.79272276E+01 1.80541406E+00 5.26493060E-02-3.30870383E-05    3
 1.04593484E-08-1.32305701E-12-1.03866773E+04 2.24829685E+01                   4
SC4H9O2                 C   4H   9O   2    0G   300.000  5000.000 1403.000     1
 1.68209433E+01 1.98834074E-02-6.71755569E-06 1.03411636E-09-5.96371075E-14    2
-1.75815350E+04-5.95731156E+01 2.27751066E+00 5.44334651E-02-3.82988187E-05    3
 1.42447767E-08-2.18864515E-12-1.25909100E+04 1.83237264E+01                   4
PC4H9O2H   8/12/15      C   4H  10O   2    0G   300.000  5000.000 1393.000     1
 1.75610913E+01 2.17832847E-02-7.46366287E-06 1.16012068E-09-6.73630029E-14    2
-3.30036118E+04-6.38547212E+01 1.04177717E+00 5.85996659E-02-3.84212378E-05    3
 1.28728231E-08-1.75491358E-12-2.70744200E+04 2.55179528E+01                   4
SC4H9O2H                C   4H  10O   2    0G   300.000  5000.000 1402.000     1
 1.78075939E+01 2.12546017E-02-7.20960281E-06 1.11291271E-09-6.43060022E-14    2
-3.48455718E+04-6.58011470E+01 1.44010868E+00 6.05300206E-02-4.36262678E-05    3
 1.66226146E-08-2.61556930E-12-2.92631492E+04 2.17354113E+01                   4
C4H8OOH1-2              C   4H   9O   2    0G   300.000  5000.000 1389.000     1
 1.67810269E+01 1.99677597E-02-6.85257220E-06 1.06628911E-09-6.19616154E-14    2
-9.14762760E+03-5.68667893E+01 2.91878364E+00 4.86143951E-02-2.81342168E-05    3
 7.64456491E-09-7.32889491E-13-3.94464787E+03 1.89326241E+01                   4
C4H8OOH1-3              C   4H   9O   2    0G   300.000  5000.000 1396.000     1
 1.61247782E+01 2.02420980E-02-6.88631475E-06 1.06534945E-09-6.16599545E-14    2
-9.16802012E+03-5.26575415E+01 2.46292502E+00 4.70131194E-02-2.42145198E-05    3
 4.65407810E-09 1.62198662E-14-3.95787917E+03 2.24569578E+01                   4
C4H8OOH1-4              C   4H   9O   2    0G   300.000  5000.000 1393.000     1
 1.69217927E+01 1.99305696E-02-6.85727522E-06 1.06879474E-09-6.21774931E-14    2
-7.87920857E+03-5.76630146E+01 1.35984095E+00 5.52812385E-02-3.75640846E-05    3
 1.32624209E-08-1.93623296E-12-2.34455867E+03 2.63197893E+01                   4
C4H8OOH2-1              C   4H   9O   2    0G   300.000  5000.000 1404.000     1
 1.77648250E+01 1.87777052E-02-6.36410476E-06 9.81958228E-10-5.67252066E-14    2
-9.93851667E+03-6.28169590E+01 2.32205003E+00 5.55032280E-02-3.97237996E-05    3
 1.47353739E-08-2.22481777E-12-4.67331585E+03 1.98332327E+01                   4
C4H8OOH2-3              C   4H   9O   2    0G   300.000  5000.000 1403.000     1
 1.70353922E+01 1.92729887E-02-6.50684653E-06 1.00126173E-09-5.77270961E-14    2
-1.09437234E+04-5.87403112E+01 3.30289851E+00 5.08231524E-02-3.39615358E-05    3
 1.17622237E-08-1.66012808E-12-6.13671017E+03 1.51726178E+01                   4
C4H8OOH2-4              C   4H   9O   2    0G   300.000  5000.000 1403.000     1
 1.72354039E+01 1.91946365E-02-6.49946502E-06 1.00210964E-09-5.78559962E-14    2
-9.71158144E+03-5.98986150E+01 1.82672511E+00 5.69912331E-02-4.24389492E-05    3
 1.67119278E-08-2.70635765E-12-4.54629884E+03 2.22051948E+01                   4
C4H8O1-2                C   4H   8O   1    0G   300.000  5000.000 1463.000     1
 1.41886108E+01 1.63162740E-02-5.16581368E-06 7.60173986E-10-4.24548403E-14    2
-2.02839382E+04-5.12817914E+01-4.29657099E+00 6.75906816E-02-5.89614134E-05    3
 2.59401158E-08-4.45926746E-12-1.48799944E+04 4.47755567E+01                   4
C4H8O1-3                C   4H   8O   1    0G   300.000  5000.000 1447.000     1
 1.32076917E+01 1.77467973E-02-5.69933762E-06 8.47771212E-10-4.77345874E-14    2
-2.11717546E+04-4.78386420E+01-5.37284363E+00 6.62224444E-02-5.35318273E-05    3
 2.19451842E-08-3.54479816E-12-1.54144887E+04 4.98345472E+01                   4
C4H8O1-4                C   4H   8O   1    0G   300.000  5000.000 1484.000     1
 1.22763349E+01 1.89105920E-02-6.09113637E-06 9.08066245E-10-5.12149503E-14    2
-2.92260872E+04-4.41235671E+01-7.78117916E+00 6.98405060E-02-5.45315920E-05    3
 2.13029617E-08-3.24666872E-12-2.28996340E+04 6.17620955E+01                   4
C4H8O2-3                C   4H   8O   1    0G   300.000  5000.000 1403.000     1
 1.06341771E+01 2.41442268E-02-1.13123977E-05 2.25480711E-09-1.54043041E-13    2
-2.10383343E+04-3.36763636E+01-4.48183187E+00 6.89313360E-02-6.15371646E-05    3
 2.73743747E-08-4.85890996E-12-1.68924193E+04 4.38882874E+01                   4
C4H8OOH1-2O2            C   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H8OOH1-3O2            C   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H8OOH1-4O2            C   4H   9O   4    0G   300.000  5000.000 1387.000     1
 2.26393370E+01 1.98017374E-02-6.92349554E-06 1.09100182E-09-6.39617643E-14    2
-2.75442161E+04-8.40747892E+01 2.91974455E+00 6.34948347E-02-4.29699499E-05    3
 1.42283155E-08-1.84506244E-12-2.04867301E+04 2.26279495E+01                   4
C4H8OOH2-1O2            C   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H8OOH2-3O2            C   4H   9O   4    0G   300.000  5000.000 1408.000     1
 2.19463055E+01 1.97307584E-02-6.65765380E-06 1.02424556E-09-5.90486257E-14    2
-3.07772334E+04-8.12053531E+01 3.34683971E+00 6.67468082E-02-5.25088611E-05    3
 2.14288389E-08-3.53381793E-12-2.47340662E+04 1.73189003E+01                   4
C4H8OOH2-4O2            C   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.15734750E+01 2.04528589E-02-6.99497777E-06 1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01 3.02241018E+00 6.53862812E-02-4.89645658E-05    3
 1.90437784E-08-3.02309317E-12-2.25805572E+04 2.05729328E+01                   4
C4H71-2,4OOH            C   4H   9O   4    0G   300.000  5000.000 1398.000     1
 2.18629952E+01 1.99359398E-02-6.85103949E-06 1.06712096E-09-6.20561893E-14    2
-2.10042547E+04-7.80706874E+01 2.99387028E+00 6.52913914E-02-4.87958562E-05    3
 1.88107554E-08-2.95256716E-12-1.46021097E+04 2.27763716E+01                   4
C4H72-1,3OOH            C   4H   9O   4    0G   300.000  5000.000 1395.000     1
 2.14626449E+01 2.02946207E-02-6.97889021E-06 1.08750673E-09-6.32605387E-14    2
-2.22196721E+04-7.60671568E+01 3.85542428E+00 6.05523559E-02-4.18122063E-05    3
 1.46680029E-08-2.07881996E-12-1.60359412E+04 1.87734959E+01                   4
C4H72-1,4OOH            C   4H   9O   4    0G   300.000  5000.000 1387.000     1
 2.10228668E+01 2.10127561E-02-7.30349553E-06 1.14623341E-09-6.70076491E-14    2
-2.02908167E+04-7.29927491E+01 3.41714555E+00 5.89885977E-02-3.76843121E-05    3
 1.18450422E-08-1.46347291E-12-1.38437952E+04 2.27094787E+01                   4
C4H71-2,3OOH            C   4H   9O   4    0G   300.000  5000.000 1406.000     1
 2.22828679E+01 1.92253507E-02-6.52860872E-06 1.00881573E-09-5.83408336E-14    2
-2.29719991E+04-8.11231836E+01 3.30790561E+00 6.66513240E-02-5.21744859E-05    3
 2.10434152E-08-3.42495389E-12-1.67536738E+04 1.95806784E+01                   4
C4H7O1-3OOH-4           C   4H   8O   3    0G   300.000  5000.000 1418.000     1
 1.87250111E+01 1.88463312E-02-6.40165949E-06 9.89754621E-10-5.72727585E-14    2
-3.29825730E+04-7.18225468E+01-5.40949665E+00 8.05102667E-02-6.64646030E-05    3
 2.73711905E-08-4.44856733E-12-2.53005240E+04 5.56327196E+01                   4
C4H7O1-3OOH-2           C   4H   8O   3    0G   300.000  5000.000 1425.000     1
 1.97110479E+01 1.79060432E-02-6.05724664E-06 9.34110479E-10-5.39628469E-14    2
-3.52532541E+04-7.83129016E+01-4.68244067E+00 8.03419743E-02-6.67264700E-05    3
 2.74081300E-08-4.41623778E-12-2.75307409E+04 5.04193128E+01                   4
C4H7O1-2OOH-4           C   4H   8O   3    0G   300.000  5000.000 1417.000     1
 1.96187267E+01 1.77382423E-02-6.03563743E-06 9.34268374E-10-5.41073277E-14    2
-3.21917914E+04-7.50295988E+01-3.06056578E+00 7.52777235E-02-6.16382083E-05    3
 2.51520765E-08-4.05109146E-12-2.49310387E+04 4.48871201E+01                   4
C4H7O1-4OOH-2           C   4H   8O   3    0G   300.000  5000.000 1470.000     1
 1.74906412E+01 1.87794733E-02-6.05491558E-06 9.03185679E-10-5.09571870E-14    2
-4.22716632E+04-6.51860330E+01-5.17426936E+00 7.89225917E-02-6.62654132E-05    3
 2.77698767E-08-4.54377840E-12-3.53780833E+04 5.35508489E+01                   4
C4H7O1-2OOH-3           C   4H   8O   3    0G   300.000  5000.000 1435.000     1
 1.83476383E+01 1.72627711E-02-5.53440131E-06 8.21396496E-10-4.61479654E-14    2
-3.29223599E+04-6.69919656E+01-9.44964311E-01 7.31026695E-02-6.71227799E-05    3
 3.12252290E-08-5.67206759E-12-2.74510619E+04 3.25427282E+01                   4
C4H7O2-3OOH-1           C   4H   8O   3    0G   300.000  5000.000 1424.000     1
 2.03028185E+01 1.69331534E-02-5.71128715E-06 8.79005552E-10-5.07088176E-14    2
-3.43451470E+04-7.95919117E+01-3.04171082E+00 7.75254740E-02-6.55776743E-05    3
 2.74944445E-08-4.52476822E-12-2.70343494E+04 4.33136810E+01                   4
C4H72-1OOH              C   4H   8O   2    0G   300.000  5000.000 1381.000     1
 1.80122740E+01 1.70340943E-02-5.89884086E-06 9.23962123E-10-5.39539803E-14    2
-1.74585465E+04-6.55209757E+01 1.29755275E+00 5.59252255E-02-4.08890003E-05    3
 1.54880526E-08-2.42412478E-12-1.16046928E+04 2.43621382E+01                   4
NC4KET12                C   4H   8O   3    0G   300.000  5000.000 1389.000     1
 2.17577434E+01 1.64473301E-02-5.79961988E-06 9.19149624E-10-5.41037382E-14    2
-4.47115295E+04-8.37725285E+01-7.24231793E-01 7.26648886E-02-6.04779190E-05    3
 2.54348857E-08-4.30152907E-12-3.72936909E+04 3.56276963E+01                   4
NC4KET13                C   4H   8O   3    0G   300.000  5000.000 1411.000     1
 1.93085398E+01 1.73455091E-02-5.85046818E-06 9.00297947E-10-5.19274609E-14    2
-4.51023813E+04-7.04869509E+01 3.31775682E+00 5.28482064E-02-3.43211665E-05    3
 1.04562704E-08-1.12796519E-12-3.94868388E+04 1.58443308E+01                   4
NC4KET14                C   4H   8O   3    0G   300.000  5000.000 1385.000     1
 1.89231898E+01 1.82270124E-02-6.27434124E-06 9.78729382E-10-5.69844333E-14    2
-4.32508875E+04-6.78717188E+01 2.92378737E+00 5.07578011E-02-2.88360718E-05    3
 6.64649914E-09-2.83907499E-13-3.72946444E+04 1.96328202E+01                   4
NC4KET21                C   4H   8O   3    0G   300.000  5000.000 1389.000     1
 2.10786402E+01 1.61788162E-02-5.53076294E-06 8.59641186E-10-4.99535144E-14    2
-4.57563821E+04-7.88014765E+01-3.88449068E-01 6.92735051E-02-5.58731127E-05    3
 2.25791086E-08-3.63900158E-12-3.86875801E+04 3.52948090E+01                   4
NC4KET23                C   4H   8O   3    0G   300.000  5000.000 1411.000     1
 1.76877593E+01 1.84820224E-02-6.18384585E-06 9.45792334E-10-5.42981801E-14    2
-4.78594254E+04-6.06681612E+01 3.56926969E+00 5.20285891E-02-3.64134216E-05    3
 1.32007682E-08-1.93576774E-12-4.30650503E+04 1.48669401E+01                   4
NC4KET24                C   4H   8O   3    0G   300.000  5000.000 1394.000     1
 1.74146206E+01 1.92744267E-02-6.57971403E-06 1.02023879E-09-5.91418353E-14    2
-4.60663138E+04-5.80320911E+01 3.12062686E+00 5.01343936E-02-3.10194950E-05    3
 9.36512355E-09-1.07548923E-12-4.08644270E+04 1.96071994E+01                   4
C4H71-3OOH              C   4H   8O   2    0G   300.000  5000.000 1392.000     1
 1.92985494E+01 1.54534427E-02-5.25460431E-06 8.13772446E-10-4.71689947E-14    2
-1.85003480E+04-7.49926639E+01-1.50977396E+00 6.85369305E-02-5.75193633E-05    3
 2.43179107E-08-4.09788488E-12-1.18018961E+04 3.50420113E+01                   4
C4H71-3,4OOH            C   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.18394783E+01 1.98802807E-02-6.81505369E-06 1.05975117E-09-6.15560073E-14    2
-2.09468667E+04-7.79984909E+01 2.56890026E+00 6.71962184E-02-5.16999792E-05    3
 2.05770379E-08-3.32914310E-12-1.45125600E+04 2.46332539E+01                   4
C4H72-3,4OOH            C   4H   9O   4    0G   300.000  5000.000 1395.000     1
 2.14626449E+01 2.02946207E-02-6.97889021E-06 1.08750673E-09-6.32605387E-14    2
-2.22196721E+04-7.60671568E+01 3.85542428E+00 6.05523559E-02-4.18122063E-05    3
 1.46680029E-08-2.07881996E-12-1.60359412E+04 1.87734959E+01                   4
HO2CH2CHO  9/ 8/14      C   2H   4O   3    0G   300.000  5000.000 1391.000     1
 1.51554685E+01 7.57240000E-03-2.72693024E-06 4.38217189E-10-2.60434287E-14    2
-3.41419680E+04-5.01255068E+01-1.32768631E+00 5.21618601E-02-4.97327645E-05    3
 2.31272366E-08-4.20787867E-12-2.90608844E+04 3.61860491E+01                   4
IC4H10     8/12/15      C   4H  10    0    0G   300.000  5000.000 1397.000     1
 1.26422737E+01 2.14133551E-02-7.26711536E-06 1.12207226E-09-6.48434177E-14    2
-2.28293782E+04-4.66059659E+01-1.07413829E+00 5.24618320E-02-3.42407949E-05    3
 1.18817533E-08-1.73238254E-12-1.79218932E+04 2.74851665E+01                   4
IC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1397.000     1
 1.23261837E+01 1.92057770E-02-6.52063623E-06 1.00704497E-09-5.82038734E-14    2
 2.50995714E+03-4.13478742E+01 1.20802408E-01 4.73187324E-02-3.16440251E-05    3
 1.14229699E-08-1.74784642E-12 6.84032915E+03 2.44291032E+01                   4
TC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1380.000     1
 1.02682832E+01 2.09965262E-02-7.14945754E-06 1.10648358E-09-6.40498314E-14    2
 1.57542675E+02-3.00960941E+01 1.05841769E+00 3.41133739E-02-9.03156779E-06    3
-2.95313136E-09 1.41436845E-12 4.22699258E+03 2.23965051E+01                   4
TC4H9O            T08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
 1.27371509E+01 2.33707342E-02-8.50516678E-06 1.38519973E-09-8.34398061E-14    2
-1.66940150E+04-4.53156321E+01 2.77057100E+00 2.68033175E-02 4.12718360E-05    3
-7.22054739E-08 3.02642276E-11-1.27079262E+04 1.21532856E+01-1.04543262E+04    4
IC4H9O            A08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
 1.16309708E+01 2.47981574E-02-9.01550536E-06 1.46714720E-09-8.83214518E-14    2
-1.37854612E+04-3.81956151E+01 3.80297372E+00 1.56874209E-02 6.81105412E-05    3
-9.83346774E-08 3.95261902E-11-1.00832243E+04 9.78963305E+00-7.82602559E+03    4
IC4H8O     9/ 1/12      C   4H   8O   1    0G   300.000  5000.000 1394.000     1
 1.40433578E+01 2.05733637E-02-9.09519220E-06 1.73417298E-09-1.14908544E-13    2
-3.62275308E+04-6.90009668E+01-5.02573822E+00 7.51340960E-02-6.88668822E-05    3
 3.12223247E-08-5.60128818E-12-3.07481413E+04 2.96284295E+01                   4
IC3H7CHO   2/22/96 THERMC   4H   8O   1    0G   300.000  5000.000 1391.000     1
 1.37501656E+01 1.83126722E-02-6.28572629E-06 9.78250756E-10-5.68538653E-14    2
-3.26936771E+04-4.77270548E+01-2.73021382E-01 4.89696307E-02-3.12770049E-05    3
 1.00052945E-08-1.27512074E-12-2.76054737E+04 2.83451139E+01                   4
IC3H7CO    2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000     1
 1.33305736E+01 1.61873930E-02-5.56711402E-06 8.67575951E-10-5.04696549E-14    2
-1.37307001E+04-4.33958746E+01 5.03452639E-01 4.41607510E-02-2.82139091E-05    3
 8.93548675E-09-1.11327422E-12-9.07755468E+03 2.61991461E+01                   4
IC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000     1
 1.33102250E+01 1.62097959E-02-5.57575891E-06 8.69003718E-10-5.05554202E-14    2
-7.62177931E+03-4.25050854E+01 5.21481767E-01 4.43114357E-02-2.86617314E-05    3
 9.30319894E-09-1.20761563E-12-2.99677086E+03 2.68182130E+01                   4
TC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1389.000     1
 1.31013047E+01 1.66391865E-02-5.68457623E-06 8.81808351E-10-5.11290161E-14    2
-1.30638647E+04-4.42705813E+01 1.87052762E+00 4.14869677E-02-2.66815701E-05    3
 9.01531610E-09-1.27870633E-12-8.97730744E+03 1.66174178E+01                   4
IC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1396.000     1
 1.33892118E+01 1.39115420E-02-4.75820958E-06 7.38736618E-10-4.28606559E-14    2
-1.97917448E+04-4.60146004E+01 1.09372823E+00 4.43315368E-02-3.41918451E-05    3
 1.39369607E-08-2.33791460E-12-1.56745978E+04 1.94458467E+01                   4
TC3H6O2CHO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1386.00      1
 1.85534443E+01 1.68774389E-02-5.90752965E-06 9.31518085E-10-5.46345187E-14    2
-2.85447191E+04-6.82486667E+01 2.17883383E+00 5.41595832E-02-3.83435886E-05    3
 1.38308104E-08-2.04190147E-12-2.27394154E+04 2.00751264E+01                   4
IC3H5O2HCHO 8/2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00      1
 2.06288832E+01 1.48625539E-02-5.25305276E-06 8.33772951E-10-4.91277401E-14    2
-2.27589076E+04-7.82962888E+01 2.05984770E+00 5.82331716E-02-4.37672100E-05    3
 1.63249918E-08-2.43462051E-12-1.63496250E+04 2.13687921E+01                   4
TC3H6O2HCO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00      1
 2.06472678E+01 1.48526500E-02-5.25104875E-06 8.33619219E-10-4.91256069E-14    2
-2.88719869E+04-7.95951389E+01 2.03864428E+00 5.80421003E-02-4.32123528E-05    3
 1.58792094E-08-2.32209543E-12-2.24284673E+04 2.03680990E+01                   4
TC3H6OCHO  8/25/95 THERMC   4H   7O   2    0G   300.000  5000.000 1394.00      1
 1.70371287E+01 1.54400645E-02-5.28332886E-06 8.21085347E-10-4.76898429E-14    2
-2.75871941E+04-6.37271230E+01 3.70830259E-01 5.38475661E-02-3.82477565E-05    3
 1.32882237E-08-1.79228730E-12-2.18391262E+04 2.58142112E+01                   4
IC3H6CO   03/03/95 THERMC   4H   6O   1    0G   300.000  5000.000 1397.00      1
 1.32548232E+01 1.40142787E-02-4.78910215E-06 7.42924342E-10-4.30737566E-14    2
-2.00529779E+04-4.44810221E+01 2.28039055E+00 4.17016989E-02-3.25089661E-05    3
 1.37243419E-08-2.40573132E-12-1.63939712E+04 1.38187714E+01                   4
IC3H5CO                 C   4H   5O   1    0G   300.000  5000.000 1396.000     1
 1.29634401E+01 1.17954996E-02-4.04361488E-06 6.28771516E-10-3.65209867E-14    2
-8.26519462E+02-4.20562575E+01 1.87306990E+00 3.95188508E-02-3.11404053E-05    3
 1.28844447E-08-2.18165308E-12 2.85270691E+03 1.68774016E+01                   4
IC3H4CHO-A              C   4H   5O   1    0G   300.000  5000.000 1392.000     1
 1.41736959E+01 1.09161978E-02-3.69020878E-06 5.69228087E-10-3.29023246E-14    2
-1.92867979E+03-5.02663740E+01 7.64345054E-01 4.45242412E-02-3.61033720E-05    3
 1.48295287E-08-2.43809290E-12 2.44732544E+03 2.08541848E+01                   4
SC4H7OH-I         L 2/00C   4H   8O   1    0G   300.000  5000.000 1395.000     1
 1.30299481E+01 1.83782479E-02-6.18529878E-06 9.49578099E-10-5.46526348E-14    2
-3.10723026E+04-4.22891828E+01 2.70103499E+00 4.17950180E-02-2.67860575E-05    3
 9.38191037E-09-1.41171285E-12-2.73561190E+04 1.35316306E+01                   4
IC4H9O2    9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1432.000     1
 1.78793870E+01 1.82474607E-02-6.01252193E-06 9.11106794E-10-5.20018932E-14    2
-1.74569774E+04-6.61552973E+01 1.77219624E+00 5.34032789E-02-3.31041810E-05    3
 9.24465657E-09-8.01706642E-13-1.17768774E+04 2.09581481E+01                   4
TC4H9O2    9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1380.000     1
 1.80863238E+01 1.99282971E-02-6.98287309E-06 1.10171726E-09-6.46381057E-14    2
-2.04420664E+04-6.97533212E+01 2.63892371E+00 5.44717499E-02-3.75504698E-05    3
 1.40479250E-08-2.27968600E-12-1.47598933E+04 1.40325533E+01                   4
IC4H8O2H-I 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1414.000     1
 1.83915486E+01 1.73042831E-02-5.66841018E-06 8.55414265E-10-4.86781778E-14    2
-9.48569748E+03-6.67673286E+01 1.86432620E-01 6.26430177E-02-4.83690886E-05    3
 1.88657148E-08-2.91189385E-12-3.59086611E+03 2.97635367E+01                   4
IC4H8O2H-T 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1413.000     1
 1.69753885E+01 1.85198010E-02-6.09075415E-06 9.21673609E-10-5.25502501E-14    2
-1.14812757E+04-5.88259039E+01 3.84374544E+00 4.36800978E-02-2.07599526E-05    3
 2.51709167E-09 5.41306513E-13-6.50766215E+03 1.34244877E+01                   4
TC4H8O2H-I 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1379.000     1
 1.81415374E+01 1.94699499E-02-6.82750014E-06 1.07773311E-09-6.32519099E-14    2
-1.23570939E+04-6.63491602E+01 3.54378349E+00 5.25201369E-02-3.69898493E-05    3
 1.44634925E-08-2.47536050E-12-6.98183185E+03 1.27623539E+01                   4
CC4H8O     9/ 1/12      C   4H   8O   1    0G   300.000  5000.000 1431.000     1
 1.51841776E+01 1.64656666E-02-5.33483091E-06 7.98149768E-10-4.51160381E-14    2
-3.33923434E+04-7.43746988E+01-6.56746688E+00 7.87298554E-02-7.33065478E-05    3
 3.40602701E-08-6.15674656E-12-2.71582518E+04 3.80875851E+01                   4
IC4H8OOH-IO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1367.000     1
 2.24664901E+01 2.09351287E-02-7.44324128E-06 1.18589255E-09-7.00546897E-14    2
-2.94495457E+04-8.54241451E+01 4.23354857E+00 5.63088857E-02-3.15672522E-05    3
 7.79536931E-09-6.21665008E-13-2.22782534E+04 1.52623111E+01                   4
IC4H8OOH-TO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1385.000     1
 2.32464612E+01 1.88384513E-02-6.40938087E-06 9.92649459E-10-5.75275879E-14    2
-3.16533132E+04-8.88301710E+01 3.36413530E+00 6.93742776E-02-5.70416393E-05    3
 2.46040165E-08-4.32848680E-12-2.51137558E+04 1.65767339E+01                   4
TC4H8OOH-IO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1385.000     1
 2.32464612E+01 1.88384513E-02-6.40938087E-06 9.92649459E-10-5.75275879E-14    2
-3.16533132E+04-8.88301710E+01 3.36413530E+00 6.93742776E-02-5.70416393E-05    3
 2.46040165E-08-4.32848680E-12-2.51137558E+04 1.65767339E+01                   4
IC4KETII   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1387.000     1
 1.95143059E+01 1.82377395E-02-6.38908606E-06 1.00801571E-09-5.91440350E-14    2
-4.46884836E+04-7.17167584E+01 1.15501614E+00 6.10622345E-02-4.49711323E-05    3
 1.70514654E-08-2.65948602E-12-3.82747956E+04 2.69612235E+01                   4
IC4KETIT   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1388.000     1
 2.09369850E+01 1.71090955E-02-6.01892169E-06 9.52353863E-10-5.59926176E-14    2
-4.77819819E+04-8.27717611E+01 1.14243741E+00 6.33840797E-02-4.73084738E-05    3
 1.77145373E-08-2.67265475E-12-4.09366796E+04 2.34844867E+01                   4
TIC4H7Q2-I 5/ 6/96 THERMC   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.33848631E+01 1.87070035E-02-6.44021945E-06 1.00428123E-09-5.84468189E-14    2
-2.61180902E+04-8.76610135E+01 4.48426361E+00 6.61225007E-02-5.27349018E-05    3
 2.18215585E-08-3.66788946E-12-1.98906586E+04 1.26719614E+01                   4
IIC4H7Q2-I 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1394.000     1
 2.30500244E+01 1.92149194E-02-6.66622576E-06 1.04495725E-09-6.10370520E-14    2
-2.32086881E+04-8.39949885E+01 4.93055661E+00 6.05819201E-02-4.23665566E-05    3
 1.49122008E-08-2.10978665E-12-1.68415495E+04 1.36228018E+01                   4
IIC4H7Q2-T 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1377.000     1
 2.15070321E+01 2.05359839E-02-7.12383399E-06 1.11655053E-09-6.52112103E-14    2
-2.51117508E+04-7.43379783E+01 8.16274487E+00 4.34463050E-02-1.76972456E-05    3
 4.88790666E-10 9.03915465E-13-1.96501749E+04 2.62067299E-01                   4
IC4H7OOH   4/15/15      C   4H   8O   2    0G   300.000  5000.000 1386.000     1
 1.82897194E+01 1.67815784E-02-5.80668193E-06 9.08949180E-10-5.30513302E-14    2
-1.82046522E+04-6.72111342E+01 1.31851762E-01 6.19561224E-02-4.99343877E-05    3
 2.09628211E-08-3.59717924E-12-1.21399925E+04 2.93905962E+01                   4
IC4H9O2H   9/ 1/12      C   4H  10O   2    0G   300.000  5000.000 1402.000     1
 1.91651624E+01 1.93678648E-02-6.41984435E-06 9.76947752E-10-5.59299558E-14    2
-3.48790978E+04-7.42063787E+01-5.47969191E-01 6.57428787E-02-4.70123149E-05    3
 1.65991096E-08-2.27331437E-12-2.82180462E+04 3.12961385E+01                   4
TC4H9O2H   9/ 1/12      C   4H  10O   2    0G   300.000  5000.000 1382.000     1
 1.90926853E+01 2.12697804E-02-7.46252626E-06 1.17841127E-09-6.91795087E-14    2
-3.77278405E+04-7.61321196E+01 4.45573540E-01 6.66153523E-02-5.20932123E-05    3
 2.22301799E-08-4.00189859E-12-3.12260714E+04 2.37278262E+01                   4
IC4H8      8/12/15      C   4H   8    0    0G   300.000  5000.000 1392.000     1
 1.11444028E+01 1.81609265E-02-6.17791116E-06 9.55481871E-10-5.52826092E-14    2
-7.84024684E+03-3.68508829E+01 5.72478139E-02 4.17768938E-02-2.49095729E-05    3
 7.54294402E-09-9.23202212E-13-3.72166259E+03 2.35698905E+01                   4
IC4H7      8/12/15      C   4H   7    0    0G   300.000  5000.000 1384.000     1
 1.18999143E+01 1.51569859E-02-5.09995449E-06 7.83722199E-10-4.51660275E-14    2
 1.00363555E+04-4.02286635E+01-2.29578762E-01 4.17842986E-02-2.66885700E-05    3
 8.42205744E-09-1.03175361E-12 1.43946680E+04 2.54797645E+01                   4
IC4H7-I1   5/13/15      C   4H   7    0    0G   300.000  5000.000 1396.000     1
 1.11158752E+01 1.55127192E-02-5.23769366E-06 8.05998394E-10-4.64703390E-14    2
 2.19488297E+04-3.41440480E+01 9.12464579E-01 3.88654394E-02-2.57575714E-05    3
 9.07760026E-09-1.33946902E-12 2.55635553E+04 2.08634918E+01                   4
IC4H7O2           L 2/00C   4H   7O   2    0G   300.000  5000.000 1404.000     1
 1.45791608E+01 1.62136068E-02-5.26957103E-06 7.90454323E-10-4.47755051E-14    2
-1.20848042E+03-4.56459433E+01 1.43532045E+00 4.89026570E-02-3.63600970E-05    3
 1.41906420E-08-2.24557878E-12 3.09284623E+03 2.41320196E+01                   4
IC4H6OOH-I        L 2/00C   4H   7O   2    0G   300.000  5000.000 1398.000     1
 1.73601429E+01 1.42046196E-02-4.65348263E-06 7.02209785E-10-3.99552775E-14    2
-1.07509366E+03-6.12822377E+01 6.06669321E+00 3.94950065E-02-2.52721718E-05    3
 7.84485641E-09-8.98876886E-13 2.87448422E+03-3.78377026E-01                   4
CCYCCOOC-T1        THERMC   4H   7O   2    0G   300.000  5000.000 1394.000     1
 1.68269657E+01 1.64471921E-02-5.63767184E-06 8.78001611E-10-5.10959632E-14    2
-3.65710841E+03-6.74096786E+01-5.29767923E+00 6.65082201E-02-4.67054235E-05    3
 1.51029775E-08-1.74322091E-12 3.97935712E+03 5.16412476E+01                   4
C2CYCOOC-I1   7/14      C   4H   7O   2    0G   300.000  5000.000 1388.000     1
 1.89745085E+01 1.50113808E-02-5.30728309E-06 8.42454740E-10-4.96392976E-14    2
-6.93111358E+03-9.08581019E+01-2.04718031E+00 7.26608379E-02-6.82960279E-05    3
 3.27505762E-08-6.23802161E-12-3.71475599E+02 1.92056057E+01                   4
IC4H7O     4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1386.000     1
 1.33457615E+01 1.61218588E-02-5.44376403E-06 8.38199374E-10-4.83608280E-14    2
 6.11443644E+02-4.36818838E+01 1.74700687E+00 4.07783436E-02-2.44750243E-05    3
 7.06502958E-09-7.51570589E-13 4.86979233E+03 1.94535999E+01                   4
CVCYCCOC          L 2/00C   4H   6O   1    0G   300.000  5000.000 1397.000     1
 1.14363523E+01 1.63250968E-02-5.57146218E-06 8.63795613E-10-5.00701899E-14    2
-5.44653450E+03-3.87179379E+01-2.45566808E+00 4.88377067E-02-3.46186324E-05    3
 1.26590643E-08-1.88737988E-12-6.43460880E+02 3.58434061E+01                   4
CCYC2OCO          L 2/00C   4H   7O   2    0G   300.000  5000.000 1401.000     1
 1.64352871E+01 1.65843210E-02-5.71790511E-06 8.92586562E-10-5.19865043E-14    2
-1.60938498E+04-5.96946106E+01-2.97381263E+00 6.75615160E-02-5.79901709E-05    3
 2.55213006E-08-4.49991674E-12-9.93607156E+03 4.25127997E+01                   4
CCYCCOOC-I2       L 2/00C   4H   7O   2    0G   300.000  5000.000 1398.000     1
 1.63388791E+01 1.65879474E-02-5.61829108E-06 8.67331033E-10-5.01476782E-14    2
 6.66946988E+03-6.40322040E+01-4.55772603E+00 7.10221387E-02-6.05228430E-05    3
 2.61773944E-08-4.51390528E-12 1.32922215E+04 4.60828737E+01                   4
CHOIC3H6O         L 2/00C   4H   7O   2    0G   300.000  5000.000 1386.000     1
 1.55511970E+01 1.67360034E-02-5.73573457E-06 8.92095191E-10-5.18351848E-14    2
-2.50674335E+04-5.23215658E+01 2.55559437E-01 5.22086026E-02-3.72283766E-05    3
 1.36714420E-08-2.05638885E-12-1.97284649E+04 2.99210251E+01                   4
IC3H5OOCH2        L 2/00C   4H   7O   2    0G   300.000  5000.000 1410.000     1
 5.05335676E+00 3.62904388E-02-1.54012992E-05 2.74341619E-09-1.74718602E-13    2
 4.08326144E+03-2.55389509E+00-1.26548168E+00-3.61337863E-03 7.31803998E-05    3
-5.49845697E-08 1.20447492E-11 1.33108969E+04 5.33428723E+01                   4
CCYCCO-T1         L 2/00C   3H   5O   1    0G   300.000  5000.000 1389.000     1
 1.03394781E+01 1.15180335E-02-3.87496644E-06 5.95744364E-10-3.43539552E-14    2
 7.17658970E+03-2.89687593E+01-1.39311392E+00 3.81789194E-02-2.62316288E-05    3
 8.74877238E-09-1.11296763E-12 1.12534953E+04 3.41877003E+01                   4
IC4H8OH-IT              C   4H   9O   1    0G   300.000  5000.000 1391.000     1
 1.29136746E+01 2.06583409E-02-6.98445966E-06 1.07562552E-09-6.20443876E-14    2
-1.81394866E+04-3.84972088E+01 3.05275715E+00 3.93926461E-02-1.90686417E-05    3
 3.86408022E-09-1.48005244E-13-1.42263749E+04 1.60840537E+01                   4
IC4H8OH-TI              C   4H   9O   1    0G   300.000  5000.000 1402.000     1
 1.46323607E+01 1.88895981E-02-6.30561450E-06 9.62474230E-10-5.51640163E-14    2
-1.87976018E+04-4.93218793E+01 2.33169342E+00 5.13017040E-02-4.02698872E-05    3
 1.75150405E-08-3.16001727E-12-1.48318978E+04 1.55368130E+01                   4
IC4H7OH                 C   4H   8O   1    0G   300.000  5000.000 1398.000     1
 1.23304221E+01 1.83885172E-02-6.06721733E-06 9.19054723E-10-5.24036171E-14    2
-2.59452023E+04-3.67418286E+01 2.04124240E+00 4.14387207E-02-2.55228632E-05    3
 8.28133017E-09-1.10654457E-12-2.22709637E+04 1.88699473E+01                   4
IC4H8OH    2/14/95 THERMC   4H   9O   1    0G   300.000  5000.000 1376.000     1
 1.25605997E+01 2.10637488E-02-7.15019648E-06 1.10439262E-09-6.38428695E-14    2
-1.86203249E+04-3.67889430E+01 3.29612707E+00 3.47649647E-02-1.02505618E-05    3
-2.04641931E-09 1.18879408E-12-1.45627247E+04 1.58606320E+01                   4
IC4H6OH                 C   4H   7O   1    0G   300.000  5000.000 1402.000     1
 1.53490714E+01 1.38856699E-02-4.56427754E-06 6.90418690E-10-3.93540403E-14    2
-1.20164758E+04-5.55975530E+01-1.46664187E+00 6.03351671E-02-5.43112644E-05    3
 2.49299933E-08-4.52282491E-12-6.95012413E+03 3.20768458E+01                   4
TQJC4H8OH               C   4H   9O   3    0G   300.000  5000.000 1415.000     1
 2.29681617E+01 1.65162786E-02-5.50247318E-06 8.39335285E-10-4.81030625E-14    2
-4.10051460E+04-9.34897892E+01-6.43419503E-01 8.49131517E-02-8.17210578E-05    3
 3.90979927E-08-7.27092842E-12-3.42375932E+04 2.84394025E+01                   4
TQC4H8OI                C   4H   9O   3    0G   300.000  5000.000 1411.000     1
 2.13200701E+01 1.80489663E-02-6.06124072E-06 9.29740751E-10-5.34977374E-14    2
-3.12966663E+04-8.20046659E+01 7.45747835E-02 7.46499596E-02-6.42255048E-05    3
 2.80908988E-08-4.87692045E-12-2.47182737E+04 2.94511549E+01                   4
QC4H7OHP                C   4H   9O   3    0G   300.000  5000.000 1416.000     1
 2.43481084E+01 1.50316366E-02-5.01788017E-06 7.66774357E-10-4.40093220E-14    2
-3.31922320E+04-9.68211106E+01-1.27864186E+00 8.94492926E-02-8.78565423E-05    3
 4.22110919E-08-7.83450876E-12-2.58975226E+04 3.53963909E+01                   4
TQC4H7OHI         L 2/00C   4H   9O   3    0G   300.000  5000.000 1404.000     1
 2.08281225E+01 1.81675094E-02-6.12943202E-06 9.43194119E-10-5.43937008E-14    2
-3.37386684E+04-7.74823720E+01 2.55843807E+00 6.37086077E-02-4.97169945E-05    3
 1.99225109E-08-3.21373436E-12-2.77526909E+04 1.95001368E+01                   4
CCY(CCO)COH             C   4H   8O   2    0G   300.000  5000.000 1412.000     1
 1.91884885E+01 1.56255714E-02-5.22569800E-06 7.99171074E-10-4.58832445E-14    2
-4.71120302E+04-7.84579023E+01-7.10048774E+00 9.53371808E-02-9.78701612E-05    3
 4.90005646E-08-9.41685766E-12-3.98987202E+04 5.60924667E+01                   4
C2CY(COC)OH             C   4H   8O   2    0G   300.000  5000.000 1393.000     1
 1.56829970E+01 1.92910506E-02-6.63718495E-06 1.03441014E-09-6.01715267E-14    2
-4.10598236E+04-5.85686221E+01 5.92324183E-01 5.52429007E-02-4.02419018E-05    3
 1.57152217E-08-2.57388393E-12-3.58241476E+04 2.23378086E+01                   4
IQJC4H8OH         L 2/00C   4H   9O   3    0G   300.000  5000.000 1410.000     1
 2.11752212E+01 1.75144254E-02-5.73227292E-06 8.63386596E-10-4.90282414E-14    2
-3.98881576E+04-8.19187015E+01 1.81448831E+00 7.47452750E-02-7.10895172E-05    3
 3.44973679E-08-6.54646593E-12-3.44023586E+04 1.77380434E+01                   4
IC3H6OHCHO              C   4H   8O   2    0G   300.000  5000.000 1393.000     1
 1.60254376E+01 1.85402212E-02-6.36973877E-06 9.91732739E-10-5.76472640E-14    2
-5.50198923E+04-5.83074874E+01 1.84080874E+00 5.29601347E-02-3.94261774E-05    3
 1.59063430E-08-2.69565279E-12-5.01437169E+04 1.75482756E+01                   4
IQC4H8OT                C   4H   9O   3    0G   300.000  5000.000 1405.000     1
 2.04823628E+01 1.82966721E-02-6.04413378E-06 9.16380548E-10-5.22866551E-14    2
-2.94287153E+04-7.53563247E+01 3.72211529E+00 6.42864861E-02-5.52809053E-05    3
 2.50036630E-08-4.53471908E-12-2.43110525E+04 1.21981167E+01                   4
IQC4H7OHT               C   4H   9O   3    0G   300.000  5000.000 1413.000     1
 2.19945886E+01 1.62011186E-02-5.23758492E-06 7.81898296E-10-4.41125515E-14    2
-3.07383725E+04-8.16613568E+01 3.58900054E+00 7.25591129E-02-7.14080484E-05    3
 3.55250907E-08-6.84991795E-12-2.57241250E+04 1.23766657E+01                   4
CCY(CCOC)OH       L 2/00C   4H   8O   2    0G   300.000  5000.000 1404.000     1
 1.43404718E+01 1.98311504E-02-6.60657660E-06 1.00779570E-09-5.77614335E-14    2
-4.30959414E+04-5.30535015E+01-2.84914896E+00 6.23736856E-02-4.70326536E-05    3
 1.84908286E-08-2.94976027E-12-3.74257004E+04 3.83163588E+01                   4
CH2COHCH2OOH            C   3H   6O   3    0G   300.000  5000.000 1398.000     1
 1.87971268E+01 1.12783442E-02-3.90789058E-06 6.12064651E-10-3.57305453E-14    2
-3.61154867E+04-6.94914300E+01-3.89823383E-01 7.01531131E-02-7.42036788E-05    3
 3.84181056E-08-7.63555985E-12-3.07879938E+04 2.86873505E+01                   4
TC3H6OH    8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000     1
 1.12222277E+01 1.36444398E-02-4.51406709E-06 7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01 1.09670360E+00 3.80727565E-02-2.75022497E-05    3
 1.07477493E-08-1.74895773E-12-1.40764487E+04 2.22475799E+01                   4
TQC4H7OHIO2             C   4H   9O   5    0G   300.000  5000.000 1402.000     1
 2.82564819E+01 1.66969871E-02-5.67314614E-06 8.78350442E-10-5.09090253E-14    2
-5.66017464E+04-1.15147927E+02 3.17336206E+00 7.94005900E-02-6.51165712E-05    3
 2.62035931E-08-4.13406290E-12-4.84943162E+04 1.77867184E+01                   4
TQC4H7OHTO2             C   4H   9O   5    0G   300.000  5000.000 1402.000     1
 2.82564819E+01 1.66969871E-02-5.67314614E-06 8.78350442E-10-5.09090253E-14    2
-5.66017464E+04-1.15147927E+02 3.17336206E+00 7.94005900E-02-6.51165712E-05    3
 2.62035931E-08-4.13406290E-12-4.84943162E+04 1.77867184E+01                   4
TQC4H7OHIQ-I            C   4H   9O   5    0G   300.000  5000.000 1384.000     1
 2.88466964E+01 1.66289773E-02-5.74301906E-06 8.98791324E-10-5.24794891E-14    2
-4.69249234E+04-1.19117836E+02 6.09881562E+00 6.93745451E-02-5.12049498E-05    3
 1.81276221E-08-2.46329781E-12-3.91393707E+04 2.93862639E+00                   4
TQC4H7OHIQ-P            C   4H   9O   5    0G   300.000  5000.000 1400.000     1
 2.81439191E+01 1.63524649E-02-5.54998081E-06 8.58603978E-10-4.97359401E-14    2
-4.84502814E+04-1.11572783E+02 3.36947511E+00 7.96855226E-02-6.74365765E-05    3
 2.82233283E-08-4.65270820E-12-4.05567534E+04 1.92726029E+01                   4
IC3H5COHQ               C   4H   8O   3    0G   300.000  5000.000 1504.000     1
 2.07387831E+01 1.58360934E-02-5.27614462E-06 8.05932218E-10-4.62682425E-14    2
-4.41821241E+04-7.94239893E+01 2.64360992E+00 5.72485066E-02-3.95907807E-05    3
 1.27775635E-08-1.47241476E-12-3.80099993E+04 1.77322273E+01                   4
CH2CQCOHQ  7/ 1/14      C   3H   6O   5    0G   300.000  5000.000 1418.000     1
 3.86574091E+01 4.83815026E-04-2.10413843E-07 3.81490832E-11-2.46187754E-15    2
-6.56392184E+04-1.61083579E+02-1.61171759E+01 1.78866440E-01-2.16751308E-04    3
 1.15450289E-07-2.27163078E-11-5.21165145E+04 1.14441286E+02                   4
IC3H5Q                  C   3H   6O   2    0G   300.000  5000.000 1397.000     1
 1.43424294E+01 1.28053632E-02-4.40584813E-06 6.86848148E-10-3.99675209E-14    2
-1.65261025E+04-4.89934539E+01 1.32903007E+00 4.49170722E-02-3.51235127E-05    3
 1.41982181E-08-2.33335008E-12-1.21898396E+04 2.02696565E+01                   4
COHQCYC(COC)            C   4H   8O   4    0G   300.000  5000.000 1319.000     1
 2.44599226E+01 1.64187782E-02-5.74024372E-06 9.05710407E-10-5.31829152E-14    2
-6.01811228E+04-1.02049722E+02 2.40687943E+00 5.95180442E-02-3.16913659E-05    3
 4.23694824E-09 8.42033474E-13-5.19694864E+04 1.88941416E+01                   4
QCYC(CCOC)OH            C   4H   8O   4    0G   300.000  5000.000 1411.000     1
 2.20860197E+01 1.83743733E-02-6.29478769E-06 9.78787994E-10-5.68621317E-14    2
-5.89652037E+04-8.64964494E+01-2.09099972E+00 8.02656739E-02-6.69756245E-05    3
 2.79282034E-08-4.60981823E-12-5.12529252E+04 4.11897260E+01                   4
HOCOCQ(CH3)2            C   4H   8O   4    0G   300.000  5000.000 1380.000     1
 2.28935401E+01 1.78627606E-02-6.34627520E-06 1.01068546E-09-5.96885712E-14    2
-8.05400680E+04-9.08953779E+01 1.56326363E+00 6.77165643E-02-5.14600149E-05    3
 1.99184629E-08-3.16007445E-12-7.30943302E+04 2.37255421E+01                   4
IQC4H7OHTO2             C   4H   9O   5    0G   300.000  5000.000 1389.000     1
 2.41720261E+01 2.09397176E-02-7.29061406E-06 1.14554056E-09-6.70217517E-14    2
-5.04772118E+04-8.95996685E+01 3.83287364E+00 6.90926177E-02-5.15031144E-05    3
 1.99235553E-08-3.17456897E-12-4.34442789E+04 1.94648622E+01                   4
IQC4H8OTQ-I             C   4H   9O   5    0G   300.000  5000.000 1386.000     1
 2.53249383E+01 2.00634820E-02-7.01249558E-06 1.10475030E-09-6.47561724E-14    2
-4.09610593E+04-9.73592779E+01 5.90219800E+00 6.26952142E-02-4.17351838E-05    3
 1.35422162E-08-1.71169663E-12-3.39620020E+04 7.89290087E+00                   4
IQC4H7OHTQ-P            C   4H   9O   5    0G   300.000  5000.000 1391.000     1
 2.45769593E+01 2.01889393E-02-7.03584537E-06 1.10623327E-09-6.47523225E-14    2
-4.25783112E+04-9.05052742E+01 3.45242802E+00 7.14541224E-02-5.54616790E-05    3
 2.22754676E-08-3.66067450E-12-3.54133076E+04 2.23024492E+01                   4
CHOC(CH3)OHCH2Q         C   4H   8O   4    0G   300.000  5000.000 1383.000     1
 2.24480753E+01 1.78753902E-02-6.26904597E-06 9.90084046E-10-5.81417382E-14    2
-6.55093075E+04-8.56747327E+01 2.40933530E+00 6.13326038E-02-4.03874986E-05    3
 1.22738404E-08-1.32997480E-12-5.83049516E+04 2.29870742E+01                   4
CO(CH2OOH)2             C   3H   6O   5    0G   300.000  5000.000 1393.000     1
 2.43376341E+01 1.14074110E-02-4.08931881E-06 6.55183244E-10-3.88570518E-14    2
-5.16862647E+04-9.01518175E+01-2.47626577E+00 8.93736793E-02-9.25891121E-05    3
 4.63168490E-08-8.93300309E-12-4.38924057E+04 4.84479477E+01                   4
CH3COCHO                C   3H   4O   2    0G   300.000  5000.000 1381.000     1
 1.14371190E+01 1.06773624E-02-3.68967757E-06 5.77006752E-10-3.36532201E-14    2
-3.78079398E+04-3.25054087E+01 2.08731049E+00 3.09032484E-02-1.98794164E-05    3
 6.26174519E-09-7.69945504E-13-3.43989451E+04 1.82839639E+01                   4
IC3H5OCH2  6/ 2/14 CZHOUH   7C   4O   1     G   298.150  2000.000 1000.00      1
 6.64731727E+00 3.08190709E-02-1.73209320E-05 5.01099629E-09-6.00089387E-13    2
 1.70679921E+03-5.91214819E+00-2.14798958E+00 7.00225553E-02-8.21595440E-05    3
 5.22589946E-08-1.34176532E-11 3.26474773E+03 3.55145589E+01                   4
IC4H7OOCH3              C   5H  10O   2    0G   300.000  5000.000 1386.000     1
 1.95896715E+01 2.31057369E-02-8.02911330E-06 1.25969946E-09-7.36169360E-14    2
-1.80069088E+04-7.34192482E+01 1.26784161E+00 6.82442475E-02-5.30807931E-05    3
 2.27496198E-08-4.11475065E-12-1.16767937E+04 2.44900544E+01                   4
IC4H7OOIC4H7            C   8H  14O   2    0G   300.000  5000.000 1390.000     1
 2.80447245E+01 3.27505220E-02-1.13220177E-05 1.77027767E-09-1.03211988E-13    2
-1.72683337E+04-1.15134796E+02-2.07881710E-01 1.04075647E-01-8.33973077E-05    3
 3.60897624E-08-6.47906520E-12-7.79062693E+03 3.50446555E+01                   4
C4H8-1                  C   4H   8    0    0G   300.000  5000.000 1388.000     1
 1.10189295E+01 1.82714177E-02-6.21801907E-06 9.62038611E-10-5.56791341E-14    2
-5.80998818E+03-3.47942287E+01 1.62599556E-01 4.01052746E-02-2.18038592E-05    3
 5.47070727E-09-4.54073315E-13-1.65402601E+03 2.48169258E+01                   4
C4H8-2     8/12/15      C   4H   8    0    0G   300.000  5000.000 1383.000     1
 1.08652083E+01 1.84123129E-02-6.26886673E-06 9.70205962E-10-5.61638967E-14    2
-7.09625867E+03-3.51547481E+01 1.30795510E+00 3.53136624E-02-1.51866126E-05    3
 1.64112363E-09 3.44257620E-13-3.19767852E+03 1.81594717E+01                   4
C4H71-1                 C   4H   7    0    0G   300.000  5000.000 1390.000     1
 1.10531750E+01 1.55668782E-02-5.25853044E-06 8.09627095E-10-4.67015477E-14    2
 2.39455759E+04-3.31548457E+01 8.97231085E-01 3.77003788E-02-2.33194855E-05    3
 7.38468124E-09-9.50027900E-13 2.76498158E+04 2.19835413E+01                   4
C4H71-2                 C   4H   7    0    0G   300.000  5000.000 1381.000     1
 1.07105686E+01 1.63539126E-02-5.63688038E-06 8.79591989E-10-5.12098725E-14    2
 2.21011255E+04-3.15300308E+01 1.56405993E+00 3.32162309E-02-1.59178310E-05    3
 2.92637814E-09-3.02645386E-14 2.57966120E+04 1.93052496E+01                   4
C4H71-3    1/13/16      C   4H   7    0    0G   300.000  5000.000 1367.000     1
 1.16977564E+01 1.53404517E-02-5.16928607E-06 7.95431212E-10-4.58914150E-14    2
 1.07395001E+04-3.82992966E+01 9.40350126E-01 3.56830321E-02-1.74384567E-05    3
 2.78964567E-09 1.78068599E-13 1.49303203E+04 2.11349333E+01                   4
C4H71-4                 C   4H   7    0    0G   300.000  5000.000 1389.000     1
 1.03875084E+01 1.63677264E-02-5.58416036E-06 8.65388736E-10-5.01415385E-14    2
 1.93282846E+04-2.86081068E+01 5.36903096E-01 3.66356251E-02-2.07814610E-05    3
 5.74895154E-09-6.05742821E-13 2.30645349E+04 2.53369983E+01                   4
C4H72-2    8/12/15      C   4H   7    0    0G   300.000  5000.000 1378.000     1
 1.05359634E+01 1.65535631E-02-5.71669066E-06 8.93155269E-10-5.20432637E-14    2
 2.08161211E+04-3.11046229E+01 2.46499885E+00 2.94957335E-02-1.08904521E-05    3
 9.17747264E-11 5.46417906E-13 2.42904093E+04 1.44728237E+01                   4
C4H71-O    4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1395.000     1
 1.53137780E+01 1.43427017E-02-4.81625517E-06 7.39574839E-10-4.26140814E-14    2
-7.29342884E+02-5.52937859E+01-1.60619192E+00 5.58562682E-02-4.35595767E-05    3
 1.70589279E-08-2.65635180E-12 4.85090326E+03 3.47112559E+01                   4
PC4H8OH-2               C   4H   9O   1    0G   300.000  5000.000 1396.000     1
 1.47198620E+01 1.93691825E-02-6.59356634E-06 1.02018538E-09-5.90410746E-14    2
-1.53023402E+04-4.85296396E+01 1.89476538E+00 4.87803114E-02-3.26702980E-05    3
 1.17119949E-08-1.77100238E-12-1.07455371E+04 2.06226225E+01                   4
SC4H8OH-1               C   4H   9O   1    0G   300.000  5000.000 1405.000     1
 1.50517242E+01 1.84748629E-02-6.15327969E-06 9.38017339E-10-5.37214281E-14    2
-1.71974443E+04-5.03733848E+01 1.78282749E+00 5.18872497E-02-3.89600849E-05    3
 1.57818686E-08-2.64133852E-12-1.28305019E+04 2.00308244E+01                   4
SC4H8OH-3               C   4H   9O   1    0G   300.000  5000.000 1403.000     1
 1.42453780E+01 1.89491000E-02-6.27403528E-06 9.52692609E-10-5.44157896E-14    2
-1.81803642E+04-4.56206494E+01 1.93185505E+00 4.79506224E-02-3.23719194E-05    3
 1.16232751E-08-1.72498918E-12-1.39431370E+04 2.03995003E+01                   4
C4H71-3OH               C   4H   8O   1    0G   300.000  5000.000 1385.000     1
 1.42401634E+01 1.83038695E-02-6.37213444E-06 1.00099740E-09-5.85511411E-14    2
-2.68183960E+04-4.83949774E+01 7.16707858E-02 5.04772909E-02-3.50356983E-05    3
 1.30539199E-08-2.07783174E-12-2.16983717E+04 2.82072724E+01                   4
C4H71-4OH               C   4H   8O   1    0G   300.000  5000.000 1396.000     1
 1.33437331E+01 1.82063693E-02-6.15150719E-06 9.47318576E-10-5.46543216E-14    2
-2.48479001E+04-4.27998774E+01-2.12276307E-01 4.86358034E-02-3.17241965E-05    3
 1.04986646E-08-1.39007078E-12-2.00365173E+04 3.04092052E+01                   4
C4H71-1OH               C   4H   8O   1    0G   300.000  5000.000 1402.000     1
 1.42586569E+01 1.71932504E-02-5.74956414E-06 8.79089774E-10-5.04586493E-14    2
-2.78051048E+04-4.96581579E+01-4.65981165E-01 5.56573217E-02-4.50578305E-05    3
 1.93726056E-08-3.38967639E-12-2.31007894E+04 2.79744544E+01                   4
C4H71-2OH               C   4H   8O   1    0G   300.000  5000.000 1404.000     1
 1.50658194E+01 1.65276030E-02-5.52197706E-06 8.43591643E-10-4.83870716E-14    2
-2.99737946E+04-5.53405024E+01-1.28560619E+00 6.35758020E-02-5.85328191E-05    3
 2.80452715E-08-5.32187122E-12-2.51538600E+04 2.93802791E+01                   4
C4H72-1OH               C   4H   8O   1    0G   300.000  5000.000 1367.000     1
 1.32893235E+01 1.93843938E-02-6.80733358E-06 1.07559847E-09-6.31698641E-14    2
-2.58627911E+04-4.34782359E+01 2.94637661E+00 3.45852975E-02-1.10024787E-05    3
-1.33281467E-09 9.54964043E-13-2.12241816E+04 1.55037145E+01                   4
C4H72-2OH               C   4H   8O   1    0G   300.000  5000.000 1402.000     1
 1.49411596E+01 1.66289929E-02-5.55627511E-06 8.48898851E-10-4.86949390E-14    2
-3.12496851E+04-5.51730870E+01-1.84033728E-01 5.90104774E-02-5.22507028E-05    3
 2.44135801E-08-4.56518659E-12-2.66717960E+04 2.36075268E+01                   4
SQC4H8OP                C   4H   9O   3    0G   300.000  5000.000 1421.000     1
 2.02482113E+01 1.90403096E-02-6.41818812E-06 9.86791658E-10-5.68666168E-14    2
-2.70686177E+04-7.43734665E+01 3.92966105E+00 5.67740736E-02-3.88077818E-05    3
 1.31554059E-08-1.72822772E-12-2.14649445E+04 1.32313419E+01                   4
PQC4H8OS                C   4H   9O   3    0G   300.000  5000.000 1403.000     1
 1.99993833E+01 1.96391125E-02-6.70755815E-06 1.04036085E-09-6.03187960E-14    2
-2.71257575E+04-7.31284601E+01 2.68979886E+00 6.10664073E-02-4.46910607E-05    3
 1.68939056E-08-2.59692346E-12-2.12460925E+04 1.94271757E+01                   4
PQC4H7OHS-3             C   4H   9O   3    0G   300.000  5000.000 1404.000     1
 1.89703648E+01 1.96512375E-02-6.61522830E-06 1.01590849E-09-5.84889733E-14    2
-2.92876345E+04-6.40682635E+01 3.14058820E+00 5.94343278E-02-4.55414505E-05    3
 1.85507067E-08-3.10109441E-12-2.40765022E+04 1.99412365E+01                   4
NC4KET12OH              C   4H   8O   2    0G   300.000  5000.000 1384.000     1
 1.68650782E+01 1.83319076E-02-6.41389893E-06 1.01105283E-09-5.92858731E-14    2
-5.27353126E+04-5.97188408E+01 5.20269850E-01 5.40316915E-02-3.57074151E-05    3
 1.18022134E-08-1.57485744E-12-4.67781081E+04 2.89999061E+01                   4
SQC4H7OHS-4             C   4H   9O   3    0G   300.000  5000.000 1414.000     1
 2.06664415E+01 1.78772156E-02-5.93193686E-06 9.02005813E-10-5.15691990E-14    2
-3.04132233E+04-7.44595459E+01 3.37952725E+00 6.50949152E-02-5.59109752E-05    3
 2.49644089E-08-4.44896795E-12-2.51501593E+04 1.58596901E+01                   4
SQC4H8OS                C   4H   9O   3    0G   300.000  5000.000 1424.000     1
 2.05363895E+01 1.85261859E-02-6.18257770E-06 9.44045247E-10-5.41390400E-14    2
-2.90453556E+04-7.66224497E+01 3.45579406E+00 6.10420456E-02-4.64106547E-05    3
 1.80687264E-08-2.81124474E-12-2.34835698E+04 1.39991890E+01                   4
NC4KET23OH    7/27/15   C   4H   8O   2    0G   300.000  5000.000 1386.000     1
 1.54636087E+01 1.92120108E-02-6.64681122E-06 1.03988604E-09-6.06552757E-14    2
-5.57292725E+04-5.19147488E+01 1.64761234E+00 4.74122084E-02-2.72508571E-05    3
 7.25755846E-09-6.68682869E-13-5.04946247E+04 2.37800424E+01                   4
SC4H8OH-3O2             C   4H   9O   3    0G   300.000  5000.000 1417.000     1
 1.93082953E+01 1.92156764E-02-6.34250732E-06 9.60912935E-10-5.47939937E-14    2
-3.84370805E+04-6.88887622E+01 1.78918281E+00 6.62988026E-02-5.52280656E-05    3
 2.40247962E-08-4.18762027E-12-3.30428157E+04 2.28885942E+01                   4
CCY(COCC)OH             C   4H   8O   2    0G   300.000  5000.000 1328.000     1
 1.03816782E+01 2.53052690E-02-1.00511826E-05 1.68204740E-09-9.58092966E-14    2
-3.94348914E+04-2.73522595E+01-6.13260697E+00 7.75376285E-02-6.73066149E-05    3
 2.82841623E-08-4.65470382E-12-3.57825027E+04 5.53089299E+01                   4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000     1
 1.12685690E+01 2.01724820E-02-7.41925667E-06 1.21275519E-09-7.30115348E-14    2
 2.13876442E+03-3.15208064E+01 5.16434924E+00 2.53427725E-02-1.39669041E-06    3
-6.00713944E-09 1.76696879E-12 5.03210693E+03 4.37441148E+00                   4
C4H6-1            L10/93C  4.H  6.   0.   0.G   200.000  6000.000 1000.        1
 7.81179394E+00 1.79733772E-02-6.61044149E-06 1.05501491E-09-6.19297169E-14    2
 1.61770171E+04-1.59658015E+01 2.42819263E+00 2.49821955E-02 6.27370548E-06    3
-2.61747866E-08 1.26585079E-11 1.80248564E+04 1.36683982E+01 1.98688798E+04    4
AC3H5OCH2  9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1397.000     1
 1.19880368E+01 1.70263516E-02-5.78617265E-06 8.94150465E-10-5.16994613E-14    2
 3.48367473E+03-3.35860630E+01 1.20089076E+00 4.24760987E-02-2.94114641E-05    3
 1.11824860E-08-1.81309530E-12 7.26792055E+03 2.43628654E+01                   4
C5H10-2    9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1385.000     1
 1.39425521E+01 2.28734997E-02-7.77800113E-06 1.20284861E-09-6.95972140E-14    2
-1.12165700E+04-4.95379542E+01 5.90528835E-01 4.85275113E-02-2.43231598E-05    3
 4.86096027E-09-1.13099201E-13-5.99777644E+03 2.41816377E+01                   4
CC5H10     9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1394.000     1
 1.44242929E+01 2.26454984E-02-7.73646334E-06 1.19999861E-09-6.95711276E-14    2
-1.14981027E+04-5.30391197E+01-9.64397004E-01 5.68482691E-02-3.66324275E-05    3
 1.23008921E-08-1.71392531E-12-5.93502026E+03 3.02998433E+01                   4
C6H10D24                C   6H  10    0    0G   300.000  5000.000 1393.000     1
 1.67662657E+01 2.32109616E-02-7.93355119E-06 1.23101995E-09-7.13892514E-14    2
-2.93324539E+03-6.44104411E+01-3.63783422E-01 6.36719104E-02-4.53090160E-05    3
 1.73368393E-08-2.79133016E-12 3.04087286E+03 2.75469470E+01                   4
C5H91-3    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1390.000     1
 1.39593933E+01 2.09180210E-02-7.14307074E-06 1.10781333E-09-6.42268160E-14    2
 7.02651017E+03-5.03103610E+01-4.68159636E-01 5.13472600E-02-3.05648794E-05    3
 8.82809744E-09-9.61458255E-13 1.23781446E+04 2.83587835E+01                   4
C5H92-4    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1384.000     1
 1.35637956E+01 2.11621316E-02-7.20826071E-06 1.11611006E-09-6.46370085E-14    2
 5.82258629E+03-4.87323606E+01 2.55028348E-01 4.69860501E-02-2.40447582E-05    3
 4.89006694E-09-1.15557679E-13 1.09775103E+04 2.46226810E+01                   4
C5H92-5    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1386.000     1
 1.32988753E+01 2.09845923E-02-7.14999241E-06 1.10717347E-09-6.41183619E-14    2
 1.39270369E+04-4.32758927E+01 9.96363945E-01 4.49148898E-02-2.30951498E-05    3
 5.01698735E-09-2.38646470E-13 1.87161506E+04 2.45616052E+01                   4
C5H91-4    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1387.000     1
 1.29229725E+01 2.10931621E-02-7.14227112E-06 1.10137556E-09-6.35983966E-14    2
 1.38192408E+04-4.00293126E+01 1.58797615E+00 4.01577239E-02-1.50062687E-05    3
-3.94608061E-10 1.02064182E-12 1.84683983E+04 2.34273438E+01                   4
C5H91-5    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1391.000     1
 1.37334869E+01 2.07003006E-02-7.06962737E-06 1.09638953E-09-6.35591113E-14    2
 1.51176253E+04-4.50794850E+01 2.07676634E-01 4.96049077E-02-3.00621602E-05    3
 9.19962077E-09-1.13246061E-12 2.01251866E+04 2.85856261E+01                   4
C5H9O2-4   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1376.000     1
 1.73707371E+01 2.09044827E-02-7.30723872E-06 1.15106814E-09-6.74601377E-14    2
-5.48020434E+03-6.50109045E+01 3.38899911E+00 4.71704753E-02-2.40389823E-05    3
 4.99166621E-09-2.03242522E-13 1.15232772E+02 1.25183625E+01                   4
SC3H5OCH2-1             C   4H   7O   1    0G   300.000  5000.000 1382.000     1
 1.47022035E+01 1.55342107E-02-5.45701052E-06 8.62544885E-10-5.06734446E-14    2
 1.81294800E+03-5.05120353E+01 2.35694446E-01 4.67367652E-02-3.04880689E-05    3
 9.75216148E-09-1.23281228E-12 7.11668364E+03 2.81378517E+01                   4
C8H141-5,3-4            C   8H  14    0    0G   300.000  5000.000 1396.000     1
 2.30690680E+01 3.23154042E-02-1.10795683E-05 1.72276354E-09-1.00052582E-13    2
-8.91240214E+03-9.49655754E+01-2.52713194E+00 9.28837673E-02-6.67176819E-05    3
 2.53683579E-08-4.01212661E-12-4.55965940E+01 4.23180878E+01                   4
C8H141-5,3  8/25/15     C   8H  14    0    0G   300.000  5000.000 1392.000     1
 2.25173982E+01 3.26748629E-02-1.11807923E-05 1.73629966E-09-1.00752481E-13    2
-8.96062790E+03-9.10857551E+01-1.02072126E+00 8.47808555E-02-5.47568199E-05    3
 1.81792070E-08-2.47335881E-12-4.53248586E+02 3.64247438E+01                   4
C8H142-6   8/25/15      C   8H  14    0    0G   300.000  5000.000 1386.000     1
 2.20960852E+01 3.27887472E-02-1.11700037E-05 1.72970378E-09-1.00179059E-13    2
-9.04951881E+03-8.92942652E+01 3.43524821E-01 7.72359120E-02-4.34861460E-05    3
 1.12949093E-08-9.77995416E-13-8.37798357E+02 2.98241439E+01                   4
C8H131-5,3-4,TA         C   8H  13    0    0G   300.000  5000.000 1394.000     1
 2.22822575E+01 3.10651867E-02-1.06940907E-05 1.66739777E-09-9.70243450E-14    2
 7.57680613E+03-9.19858764E+01-3.23996819E+00 9.13494930E-02-6.60037456E-05    3
 2.51706078E-08-3.99030974E-12 1.64345368E+04 4.49498860E+01                   4
C8H131-5,3,TA           C   8H  13    0    0G   300.000  5000.000 1389.000     1
 2.16161787E+01 3.14326704E-02-1.07786324E-05 1.67632587E-09-9.73755313E-14    2
 7.60897211E+03-8.80384104E+01-5.03201172E-01 7.78854227E-02-4.63156182E-05    3
 1.32834166E-08-1.42623050E-12 1.58388712E+04 3.26514434E+01                   4
C8H131-5,3,SA           C   8H  13    0    0G   300.000  5000.000 1392.000     1
 2.21141889E+01 3.09871348E-02-1.06198459E-05 1.65100088E-09-9.58788408E-14    2
 8.08509780E+03-9.01448021E+01-1.32185914E+00 8.30473789E-02-5.42213233E-05    3
 1.80737386E-08-2.45105483E-12 1.65183103E+04 3.67169651E+01                   4
C8H131-5,3,PA           C   8H  13    0    0G   300.000  5000.000 1389.000     1
 2.32085707E+01 2.97529224E-02-1.01333635E-05 1.56925634E-09-9.09001242E-14    2
 8.95338901E+03-9.40777602E+01-1.57063382E+00 8.60080913E-02-5.83884368E-05    3
 2.02048105E-08-2.83115953E-12 1.77015232E+04 3.95476224E+01                   4
C8H132-6,SA             C   8H  13    0    0G   300.000  5000.000 1387.000     1
 2.16167233E+01 3.12260643E-02-1.06640216E-05 1.65409816E-09-9.59112187E-14    2
 8.03384556E+03-8.72194430E+01 2.20017932E-01 7.48621425E-02-4.21239973E-05    3
 1.07414215E-08-8.66560315E-13 1.61027987E+04 2.99517204E+01                   4
C8H132-6,PA             C   8H  13    0    0G   300.000  5000.000 1378.000     1
 2.29293875E+01 2.97187394E-02-1.00712335E-05 1.55505094E-09-8.99129602E-14    2
 8.77975921E+03-9.24517461E+01 1.05119796E-01 7.70150350E-02-4.48890925E-05    3
 1.19516688E-08-1.04377517E-12 1.72713386E+04 3.22058738E+01                   4
C6H101-3,3              C   6H  10    0    0G   300.000  5000.000 1395.000     1
 1.69678361E+01 2.28868236E-02-7.78758381E-06 1.20465198E-09-6.97080856E-14    2
-2.97276905E+03-6.58632941E+01-3.01310455E-02 6.43105079E-02-4.75083462E-05    3
 1.89877768E-08-3.17681035E-12 2.82367411E+03 2.49254708E+01                   4
C8H131-5,3-4,TAO        C   8H  13O   1    0G   300.000  5000.000 1394.000     1
 2.70579050E+01 2.84726632E-02-9.66434779E-06 1.49337149E-09-8.63788413E-14    2
-4.43111126E+03-1.12228392E+02 1.00679908E+00 8.90191278E-02-6.27963646E-05    3
 2.24161585E-08-3.20587060E-12 4.56422741E+03 2.76546640E+01                   4
C8H131-5,3,TAO          C   8H  13O   1    0G   300.000  5000.000 1396.000     1
 2.16638860E+01 2.77253448E-02-9.69375951E-06 1.67582120E-09-1.08059396E-13    2
-5.70300683E+03-9.33237797E+01 1.46771925E+00 7.67800622E-02-5.63189881E-05    3
 2.22689786E-08-3.64813515E-12 1.17475936E+03 1.45619856E+01                   4
C8H131-5,3,SAO          C   8H  13O   1    0G   300.000  5000.000 1385.000     1
 2.61023602E+01 3.05036647E-02-1.06268215E-05 1.67026867E-09-9.77389024E-14    2
-3.64744193E+03-1.06781316E+02 1.60953926E+00 8.39738786E-02-5.49469234E-05    3
 1.84255257E-08-2.56040058E-12 5.33713436E+03 2.62653941E+01                   4
C8H131-5,3,PAO          C   8H  13O   1    0G   300.000  5000.000 1374.000     1
 2.51902631E+01 3.15630048E-02-1.10568300E-05 1.74424175E-09-1.02327221E-13    2
-1.34401684E+03-1.01448477E+02 3.91532442E+00 7.10319966E-02-3.55623644E-05    3
 6.98595095E-09-1.83465840E-13 7.22911524E+03 1.67145758E+01                   4
C8H132-6,SAO            C   8H  13O   1    0G   300.000  5000.000 1381.000     1
 2.54267504E+01 3.10421548E-02-1.08045689E-05 1.69716523E-09-9.92701997E-14    2
-3.28641768E+03-1.02872762E+02 3.34168622E+00 7.49917518E-02-4.18382842E-05    3
 1.06108028E-08-8.96488454E-13 5.24458399E+03 1.86128166E+01                   4
C8H132-6,PAO            C   8H  13O   1    0G   300.000  5000.000 2014.000     1
 1.99391776E+01 3.79081645E-02-1.37893231E-05 2.23770591E-09-1.34044177E-13    2
 1.42981257E+03-7.07923233E+01 6.30807632E+00 5.80374259E-02-1.75637726E-05    3
-2.70887760E-09 1.61702129E-12 7.07839485E+03 6.29344560E+00                   4
C7H111-5,3,6P           C   7H  11    0    0G   300.000  5000.000 1396.000     1
 1.95787047E+01 2.54213538E-02-8.68127275E-06 1.34629701E-09-7.80464853E-14    2
 2.58537943E+04-7.44112330E+01-6.76848821E-01 7.38082653E-02-5.35945220E-05    3
 2.06293915E-08-3.29701110E-12 3.28160434E+04 3.40518079E+01                   4
C7H111-5,1P             C   7H  11    0    0G   300.000  5000.000 1388.000     1
 1.91915682E+01 2.55013021E-02-8.65881522E-06 1.33796943E-09-7.73784878E-14    2
 2.60946287E+04-7.21387547E+01 8.16831855E-01 6.56745024E-02-4.14490949E-05    3
 1.32234876E-08-1.69289568E-12 3.27646149E+04 2.75442934E+01                   4
C4H64,2-1OH             C   4H   7O   1    0G   300.000  5000.000 1366.000     1
 1.36259446E+01 1.70233137E-02-6.00460246E-06 9.51603754E-10-5.60055773E-14    2
-7.81498890E+03-4.44948073E+01 2.50804582E+00 3.53393033E-02-1.41418095E-05    3
 5.65501810E-10 5.94838384E-13-3.08574102E+03 1.81061546E+01                   4
C4H63,1-1OH             C   4H   7O   1    0G   300.000  5000.000 1401.000     1
 1.38675222E+01 1.54795810E-02-5.17720236E-06 7.91828077E-10-4.54656891E-14    2
-1.07655481E+04-4.87820652E+01-5.96640682E-01 5.31885124E-02-4.34791765E-05    3
 1.86514084E-08-3.23780972E-12-6.15543596E+03 2.74734171E+01                   4
C4H63,1-3OH             C   4H   7O   1    0G   300.000  5000.000 1380.000     1
 1.33633351E+01 1.70222596E-02-5.95245190E-06 9.37896168E-10-5.49767305E-14    2
-9.90113178E+03-4.54753472E+01 5.96155469E-01 4.35893351E-02-2.65985265E-05    3
 8.14250262E-09-1.02316366E-12-5.05630797E+03 2.43923636E+01                   4
C4H63,1-2OH             C   4H   7O   1    0G   300.000  5000.000 1404.000     1
 1.46899596E+01 1.48008021E-02-4.94483770E-06 7.55542892E-10-4.33461574E-14    2
-1.29448240E+04-5.45653093E+01-1.58903600E+00 6.17722944E-02-5.78263835E-05    3
 2.78090017E-08-5.26779799E-12-8.17977186E+03 2.96999338E+01                   4
C4H5OH-13  9/24/15      C   4H   6O   1    0G   300.000  5000.000 1405.000     1
 1.40975061E+01 1.29826578E-02-4.36356696E-06 6.69260196E-10-3.84920001E-14    2
-1.41099189E+04-4.94340793E+01-1.60022758E+00 6.12386329E-02-6.18933585E-05    3
 3.14927455E-08-6.20396658E-12-9.77435172E+03 3.08328186E+01                   4
SQC4H7OHP-4             C   4H   9O   3    0G   300.000  5000.000 1410.000     1
 1.99207495E+01 1.89422879E-02-6.39488327E-06 9.84231371E-10-5.67606301E-14    2
-2.89250584E+04-7.01061222E+01 1.44518283E+00 6.52944119E-02-5.10380130E-05    3
 2.05238910E-08-3.32050656E-12-2.29059890E+04 2.78546218E+01                   4
CY(CCCO)COH             C   4H   8O   2    0G   300.000  5000.000 1396.000     1
 1.34636332E+01 2.28745777E-02-9.93619553E-06 1.89605197E-09-1.26466856E-13    2
-3.96396606E+04-4.51064489E+01-6.97589766E+00 7.98392838E-02-7.11131714E-05    3
 3.16611877E-08-5.61324136E-12-3.35777839E+04 6.12093340E+01                   4
NC4KET21OH              C   4H   8O   2    0G   300.000  5000.000 1507.000     1
 1.52252911E+01 1.86615017E-02-6.30658772E-06 9.72355897E-10-5.61770184E-14    2
-5.34759661E+04-5.00397269E+01 5.46677192E+00 3.01119974E-02-2.59548850E-06    3
-7.61700554E-09 2.55573161E-12-4.89909104E+04 6.33307684E+00                   4
C2H5CHOHCO              C   4H   7O   2    0G   300.000  5000.000 1389.000     1
 1.82917246E+01 1.48007410E-02-5.24974573E-06 8.35220286E-10-4.92942253E-14    2
-3.36703722E+04-7.12363783E+01-2.44749259E+00 6.46308488E-02-5.10457937E-05    3
 1.99850773E-08-3.12214490E-12-2.66670442E+04 3.95566556E+01                   4
CH3COCOHCH3             C   4H   7O   2    0G   300.000  5000.000 1395.000     1
 1.65624631E+01 1.59037217E-02-5.54554278E-06 8.72274939E-10-5.10735025E-14    2
-3.65884887E+04-6.10833920E+01-1.65607674E+00 6.08409982E-02-4.85215440E-05    3
 1.97794382E-08-3.26305133E-12-3.05158227E+04 3.58911868E+01                   4
C2H4COCH2OH             C   4H   7O   2    0G   300.000  5000.000 1462.000     1
 1.40828195E+01 1.76833414E-02-6.09759192E-06 9.52794521E-10-5.55571628E-14    2
-3.37518398E+04-4.08944306E+01 7.98874348E+00 1.41152447E-02 1.86299924E-05    3
-1.99223089E-08 5.12983835E-12-2.98706372E+04-1.87192030E+00                   4
CH3COHCO   9/24/15      C   3H   4O   2    0G   300.000  5000.000 1410.000     1
 1.50110709E+01 7.26697312E-03-2.42872486E-06 3.71246886E-10-2.13068531E-14    2
-3.87354954E+04-5.41005540E+01 8.25855205E-01 5.22217422E-02-5.66992291E-05    3
 2.94815948E-08-5.81714952E-12-3.50157127E+04 1.78488731E+01                   4
CH2COHCHO  9/24/15      C   3H   4O   2    0G   300.000  5000.000 1406.000     1
 1.40200417E+01 7.95092924E-03-2.63244516E-06 3.99896432E-10-2.28538120E-14    2
-3.76808145E+04-4.80457990E+01 5.76639663E-02 5.16589617E-02-5.49773816E-05    3
 2.83487148E-08-5.57464421E-12-3.39594513E+04 2.29757289E+01                   4
SQC4H7OHP-4O2           C   4H   9O   5    0G   300.000  5000.000 1402.000     1
 2.35936348E+01 2.08588461E-02-7.13602285E-06 1.10820581E-09-6.43133049E-14    2
-4.78452356E+04-8.49505816E+01 2.62618431E+00 7.26812595E-02-5.64956508E-05    3
 2.25892409E-08-3.65246549E-12-4.08999596E+04 2.65615323E+01                   4
PQC4H7OHS-3O2           C   4H   9O   5    0G   300.000  5000.000 1414.000     1
 2.46607662E+01 1.92947770E-02-6.45433722E-06 9.87246207E-10-5.66889630E-14    2
-4.98467067E+04-9.10424907E+01 2.90986916E+00 7.76596028E-02-6.68513896E-05    3
 2.93627835E-08-5.12008013E-12-4.31551961E+04 2.29130715E+01                   4
SQC4H7OHS-4O2           C   4H   9O   5    0G   300.000  5000.000 1414.000     1
 2.46607662E+01 1.92947770E-02-6.45433722E-06 9.87246207E-10-5.66889630E-14    2
-4.98467067E+04-9.10424907E+01 2.90986916E+00 7.76596028E-02-6.68513896E-05    3
 2.93627835E-08-5.12008013E-12-4.31551961E+04 2.29130715E+01                   4
C4H7O2-1,3OOH           C   4H   9O   5    0G   300.000  5000.000 1425.000     1
 2.54691227E+01 1.86441036E-02-6.23825706E-06 9.54422873E-10-5.48154425E-14    2
-4.01531561E+04-9.60389710E+01 4.88339443E+00 7.18219147E-02-5.86792171E-05    3
 2.42823866E-08-3.98538527E-12-3.36575518E+04 1.24696185E+01                   4
NC4KET13OH-2            C   4H   8O   4    0G   300.000  5000.000 1395.000     1
 2.25434165E+01 1.76377030E-02-6.14926113E-06 9.67201484E-10-5.66321794E-14    2
-6.59724022E+04-8.48522697E+01 2.13332105E+00 6.69840817E-02-5.19672275E-05    3
 2.03864253E-08-3.22074763E-12-5.90962942E+04 2.40964870E+01                   4
NC4KET24OH-1            C   4H   8O   4    0G   300.000  5000.000 1672.000     1
 1.76639507E+01 2.38921914E-02-8.87612081E-06 1.46065294E-09-8.83476797E-14    2
-6.36561283E+04-5.60405234E+01 7.17383002E+00 3.72830917E-02-7.30000099E-06    3
-5.42423663E-09 1.94298976E-12-5.91469605E+04 3.98040888E+00                   4
NC4KET24OH-3            C   4H   8O   4    0G   300.000  5000.000 1392.000     1
 2.02237496E+01 1.94540798E-02-6.73928381E-06 1.05529414E-09-6.15931037E-14    2
-6.68651215E+04-6.99676945E+01 2.60979522E+00 6.11530456E-02-4.50409252E-05    3
 1.73313054E-08-2.75573967E-12-6.07708447E+04 2.44892030E+01                   4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000     1
 2.15163584E+01 1.55811846E-02-5.27569793E-06 8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00 7.72727339E-02-6.79667571E-05    3
 2.98158102E-08-5.16343458E-12-3.01649655E+04 4.06810164E+01                   4
C4H6OHOOH2-2-1          C   4H   8O   3    0G   300.000  5000.000 1396.000     1
 2.16656460E+01 1.59965487E-02-5.52214578E-06 8.62740322E-10-5.02768063E-14    2
-4.14875437E+04-8.39377540E+01 4.72576793E-02 7.85787048E-02-7.68006410E-05    3
 3.79206120E-08-7.33203833E-12-3.51140091E+04 2.80064858E+01                   4
C4H6OHOOH1-3-4          C   4H   8O   3    0G   300.000  5000.000 1391.000     1
 1.93445152E+01 1.82185729E-02-6.34491630E-06 9.97097673E-10-5.83420009E-14    2
-3.79952136E+04-6.88144861E+01 9.44277749E-01 6.34330602E-02-4.99455695E-05    3
 2.05720571E-08-3.48143957E-12-3.17827282E+04 2.92923796E+01                   4
C4H6OHOOH1-2-3          C   4H   8O   3    0G   300.000  5000.000 1403.000     1
 2.32793098E+01 1.38280934E-02-4.61330737E-06 7.05319574E-10-4.05174739E-14    2
-4.26348237E+04-9.51979841E+01-2.88475927E+00 9.16099207E-02-9.37152074E-05    3
 4.66406895E-08-8.92736049E-12-3.52899912E+04 3.92851633E+01                   4
HOCH2CHO   9/24/15      C   2H   4O   2    0G   300.000  5000.000 1680.000     1
 7.99598542E+00 1.20664034E-02-4.43693399E-06 7.25167046E-10-4.36535460E-14    2
-4.09020567E+04-1.33754312E+01 4.35084369E+00 1.50412895E-02-5.95083030E-07    3
-3.75736217E-09 1.09353598E-12-3.91654526E+04 8.09610238E+00                   4
C4H71-4OOH              C   4H   8O   2    0G   300.000  5000.000 1392.000     1
 1.59871304E+01 1.86028119E-02-6.40003189E-06 9.97531711E-10-5.80334203E-14    2
-1.70152141E+04-5.46227137E+01 1.31653247E+00 5.16546159E-02-3.47310922E-05    3
 1.20405755E-08-1.71650639E-12-1.17754576E+04 2.46384545E+01                   4
C4H71-4O2  9/25/15      C   4H   7O   2    0G   300.000  5000.000 1390.000     1
 1.50240251E+01 1.72860962E-02-5.94297061E-06 9.25861430E-10-5.38461748E-14    2
 1.92460667E+02-4.85941022E+01 2.09042625E+00 4.57130080E-02-2.94815830E-05    3
 9.69604853E-09-1.30061388E-12 4.88932667E+03 2.15456077E+01                   4
C4H61-3OOH4             C   4H   7O   2    0G   300.000  5000.000 1391.000     1
 1.55818475E+01 1.69176098E-02-5.84009100E-06 9.12401042E-10-5.31699330E-14    2
 1.20753065E+01-5.36683745E+01 1.00320366E+00 4.99893791E-02-3.43100656E-05    3
 1.20104294E-08-1.71132691E-12 5.17744264E+03 2.49842453E+01                   4
C4H6O1-3OOH4            C   4H   7O   3    0G   300.000  5000.000 1386.000     1
 1.95456291E+01 1.60358540E-02-5.61768950E-06 8.86341914E-10-5.20072732E-14    2
-1.12679434E+04-6.99490153E+01 3.83045773E+00 5.07388403E-02-3.42226447E-05    3
 1.13486298E-08-1.48529245E-12-5.61786232E+03 1.51509867E+01                   4
C4H6O2-1OOH4            C   4H   7O   3    0G   300.000  5000.000 1364.000     1
 2.05164800E+01 1.55727845E-02-5.54197222E-06 8.83592649E-10-5.22241946E-14    2
-9.30030707E+03-7.46630628E+01 5.38344712E+00 4.47089832E-02-2.43630482E-05    3
 5.07835349E-09-1.20805939E-13-3.40711224E+03 8.84731441E+00                   4
HOCH2COCH2              C   3H   5O   2    0G   300.000  5000.000 1363.000     1
 1.27106963E+01 1.15513960E-02-3.95951917E-06 6.16237371E-10-3.58328248E-14    2
-2.71538154E+04-3.67129478E+01 4.98634970E+00 2.51766916E-02-1.10893306E-05    3
 1.12011467E-09 2.89491135E-13-2.40047973E+04 6.38258616E+00                   4
HOCH2CO    9/25/15      C   2H   3O   2    0G   300.000  5000.000 1487.000     1
 9.43496508E+00 7.68897340E-03-2.74959280E-06 4.39772312E-10-2.60488233E-14    2
-2.29700136E+04-2.04618579E+01 5.12916864E+00 9.07172819E-03 6.49228146E-06    3
-8.56591893E-09 2.31070825E-12-2.06151607E+04 5.73007596E+00                   4
HOCHCHO    9/25/15      C   2H   3O   2    0G   300.000  5000.000 1680.000     1
 9.99251726E+00 7.77560619E-03-2.94238616E-06 4.90136333E-10-2.98979778E-14    2
-2.20440827E+04-2.73957153E+01 5.42856274E-01 2.95295948E-02-2.08315490E-05    3
 6.72777461E-09-8.06116446E-13-1.89378452E+04 2.31681075E+01                   4
PC3H4OH-3  9/25/15      C   3H   5O   1    0G   300.000  5000.000 1378.000     1
 1.15297558E+01 1.14381097E-02-4.04415495E-06 6.41949269E-10-3.78242456E-14    2
-3.45486444E+03-3.65385497E+01 4.06368169E-01 3.70231405E-02-2.72202689E-05    3
 1.05783475E-08-1.73632514E-12 5.27160824E+02 2.34781848E+01                   4
PC3H4OH-1  9/25/15      C   3H   5O   1    0G   300.000  5000.000 1403.000     1
 1.09468986E+01 1.04014540E-02-3.44082448E-06 5.22105632E-10-2.98049266E-14    2
 4.11530600E+03-3.11161699E+01 2.07150195E+00 3.50016810E-02-3.01922013E-05    3
 1.38467853E-08-2.55380109E-12 6.81914209E+03 1.51916605E+01                   4
CH3COCHOH  9/25/15      C   3H   5O   2    0G   300.000  5000.000 1378.000     1
 1.23884831E+01 1.23099892E-02-4.32263800E-06 6.83043939E-10-4.01192794E-14    2
-2.97609476E+04-3.85682589E+01 2.11183979E+00 3.32521318E-02-1.96834015E-05    3
 5.40736760E-09-5.32450556E-13-2.58545486E+04 1.77643465E+01                   4
SC2H2OH    9/25/15      C   2H   3O   1    0G   300.000  5000.000 1410.000     1
 7.99235139E+00 5.83109353E-03-1.89242965E-06 2.83129118E-10-1.59933287E-14    2
 9.51237374E+03-1.62058375E+01 1.63791895E+00 2.64968839E-02-2.74821415E-05    3
 1.43110557E-08-2.85794966E-12 1.11467016E+04 1.58714777E+01                   4
PC4H8OH-1               C   4H   9O   1    0G   300.000  5000.000 1392.000     1
 1.47813217E+01 1.89692972E-02-6.38671427E-06 9.81341181E-10-5.65332084E-14    2
-1.88487062E+04-4.98892364E+01 7.72566991E-01 5.00429367E-02-3.20163534E-05    3
 1.02913291E-08-1.30709217E-12-1.38421800E+04 2.58928300E+01                   4
PC4H8OH-3               C   4H   9O   1    0G   300.000  5000.000 1398.000     1
 1.45944628E+01 1.92223378E-02-6.48868808E-06 9.98309067E-10-5.75488987E-14    2
-1.52392636E+04-4.85127747E+01 2.21685429E+00 4.71340178E-02-3.04254756E-05    3
 1.03165429E-08-1.45043599E-12-1.08208508E+04 1.83497891E+01                   4
C4H7O1-4   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1388.000     1
 1.33251126E+01 1.65057558E-02-5.65235890E-06 8.78319847E-10-5.09914580E-14    2
 1.91281414E+03-4.28181479E+01 2.44895430E+00 3.69423519E-02-1.77510852E-05    3
 2.64537530E-09 2.43666218E-13 6.16385921E+03 1.73174889E+01                   4
PC4H8OH-4               C   4H   9O   1    0G   300.000  5000.000 1401.000     1
 1.41519859E+01 1.96439700E-02-6.64537615E-06 1.02402720E-09-5.91001981E-14    2
-1.56141213E+04-4.50604102E+01-6.95634735E-02 5.20263179E-02-3.44849029E-05    3
 1.17704221E-08-1.63047436E-12-1.06053581E+04 3.15909567E+01                   4
SC4H8OH-2               C   4H   9O   1    0G   300.000  5000.000 1395.000     1
 1.45514712E+01 1.92722299E-02-6.50955109E-06 1.00200009E-09-5.77830714E-14    2
-2.09909632E+04-4.82454428E+01 1.96361387E+00 4.77673982E-02-3.11652479E-05    3
 1.07498897E-08-1.54834306E-12-1.65000330E+04 1.97286755E+01                   4
CH2COHCO   9/25/15      C   3H   3O   2    0G   300.000  5000.000 1411.000     1
 1.31285142E+01 6.17948608E-03-1.93387986E-06 2.81892606E-10-1.56244314E-14    2
-1.93507932E+04-4.22958094E+01 1.24341370E+00 4.71484739E-02-5.44200189E-05    3
 2.95970356E-08-6.01447282E-12-1.65555219E+04 1.68301276E+01                   4
C4H72-2O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1390.000     1
 1.63301022E+01 1.60698895E-02-5.50238293E-06 8.55098973E-10-4.96517196E-14    2
-4.70039715E+03-5.78736400E+01 2.49537080E+00 4.75680882E-02-3.26452548E-05    3
 1.14069694E-08-1.61494862E-12 1.76383849E+02 1.67027189E+01                   4
C4H71-1O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1390.000     1
 1.63738534E+01 1.62685376E-02-5.62192103E-06 8.78982520E-10-5.12510706E-14    2
-1.06318473E+03-5.69005716E+01 2.02223104E+00 4.85577506E-02-3.30293697E-05    3
 1.13406677E-08-1.57078109E-12 4.04143594E+03 2.06106646E+01                   4
C4H71-2O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1394.000     1
 1.63565639E+01 1.61768136E-02-5.56610316E-06 8.67700997E-10-5.04886444E-14    2
-3.40245466E+03-5.75260769E+01 1.42459973E+00 5.20547601E-02-3.89440869E-05    3
 1.51726193E-08-2.42611664E-12 1.68854104E+03 2.23230947E+01                   4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000     1
 1.14795375E+01 1.45881429E-02-4.88359380E-06 7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01 1.13614529E+00 3.68850655E-02-2.24073579E-05    3
 6.62398992E-09-7.32206246E-13-1.09273174E+04 2.24919343E+01                   4
PC4H8OH-2O2             C   4H   9O   3    0G   300.000  5000.000 1407.000     1
 1.90513685E+01 2.00624257E-02-6.76970282E-06 1.04136985E-09-6.00271674E-14    2
-3.65966815E+04-6.71202048E+01 1.97780900E+00 6.25692373E-02-4.76730210E-05    3
 1.90561997E-08-3.10596799E-12-3.09625439E+04 2.35880251E+01                   4
SC4H8OH-1O2             C   4H   9O   3    0G   300.000  5000.000 1405.000     1
 1.88547090E+01 2.02217653E-02-6.82328766E-06 1.04961552E-09-6.05032676E-14    2
-3.65721162E+04-6.59105449E+01 1.47037864E+00 6.38295256E-02-4.92333916E-05    3
 1.99704964E-08-3.30499356E-12-3.08602292E+04 2.63462505E+01                   4
C4H71-3OOCH3            C   5H  10O   2    0G   300.000  5000.000 1387.000     1
 2.12299326E+01 2.07003584E-02-6.99464238E-06 1.07836941E-09-6.22999849E-14    2
-1.85005682E+04-8.53499854E+01-5.42404662E-01 7.51511469E-02-6.00684679E-05    3
 2.49701271E-08-4.22319878E-12-1.13061371E+04 3.02981962E+01                   4
C4H72-1OOCH3            C   5H  10O   2    0G   300.000  5000.000 1382.000     1
 1.92914755E+01 2.34475159E-02-8.16713690E-06 1.28338262E-09-7.50837828E-14    2
-1.72688938E+04-7.16509708E+01 2.44675386E+00 6.21430218E-02-4.39326296E-05    3
 1.72567499E-08-2.94950711E-12-1.11431755E+04 1.94028997E+01                   4
C4H6                    C   4H   6    0    0G   300.000  5000.000 1388.000     1
 1.01064561E+01 1.46248415E-02-5.01373934E-06 7.79510645E-10-4.52675769E-14    2
 9.96133753E+03-2.97310638E+01 1.01356056E+00 3.35722771E-02-1.96279376E-05    3
 5.74803850E-09-6.75029065E-13 1.33956759E+04 1.99957382E+01                   4
C4H612            A 8/83C   4H   6    0    0G   300.000  5000.000 1374.000     1
 1.14059885E+01 1.31489843E-02-4.43542071E-06 6.83028825E-10-3.94289265E-14    2
 1.42427294E+04-3.69674067E+01 9.45515689E-01 3.46162239E-02-1.98590697E-05    3
 5.02139421E-09-3.67977164E-13 1.81439079E+04 2.02191143E+01                   4
C4H6-2            A 8/83C   4H   6    0    0G   300.000  5000.000 1377.000     1
 9.60305554E+00 1.48972169E-02-5.16751230E-06 8.09757170E-10-4.72817668E-14    2
 1.24831314E+04-2.87129792E+01 1.97152408E+00 2.76790997E-02-1.13396645E-05    3
 1.02970745E-09 2.75290944E-13 1.57283766E+04 1.42147356E+01                   4
C4H5-I            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 0.10229092E+02 0.94850138E-02-0.90406445E-07-0.12596100E-08 0.24781468E-12    2
 0.34642812E+05-0.28564529E+02-0.19932900E-01 0.38005672E-01-0.27559450E-04    3
 0.77835551E-08 0.40209383E-12 0.37496223E+05 0.24394241E+02                   4
C4H5-N            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 0.98501978E+01 0.10779008E-01-0.13672125E-05-0.77200535E-09 0.18366314E-12    2
 0.38840301E+05-0.26001846E+02 0.16305321E+00 0.39830137E-01-0.34000128E-04    3
 0.15147233E-07-0.24665825E-11 0.41429766E+05 0.23536163E+02                   4
C4H5-2            H6W/94C   4H   5    0    0G   300.000  5000.000 1385.000     1
 1.03230828E+01 1.17625574E-02-4.00004665E-06 6.18727929E-10-3.58083530E-14    2
 3.25861413E+04-2.88794317E+01 2.31011292E+00 2.83747046E-02-1.63836755E-05    3
 4.46251967E-09-4.30510879E-13 3.55842945E+04 1.49105965E+01                   4
C4H4              H6W/94C   4H   4    0    0G   300.000  3000.00  1000.00      1
 0.66507092E+01 0.16129434E-01-0.71938875E-05 0.14981787E-08-0.11864110E-12    2
 0.31195992E+05-0.97952118E+01-0.19152479E+01 0.52750878E-01-0.71655944E-04    3
 0.55072423E-07-0.17286228E-10 0.32978504E+05 0.31419983E+02                   4
C4H3-I            AB1/93C   4H   3    0    0G   300.000  3000.00  1000.00      1
 0.90978165E+01 0.92207119E-02-0.33878441E-05 0.49160498E-09-0.14529780E-13    2
 0.56600574E+05-0.19802597E+02 0.20830412E+01 0.40834274E-01-0.62159685E-04    3
 0.51679358E-07-0.17029184E-10 0.58005129E+05 0.13617462E+02                   4
C4H3-N            H6W/94C   4H   3    0    0G   300.000  3000.00  1000.00      1
 0.54328279E+01 0.16860981E-01-0.94313109E-05 0.25703895E-08-0.27456309E-12    2
 0.61600680E+05-0.15673981E+01-0.31684113E+00 0.46912100E-01-0.68093810E-04    3
 0.53179921E-07-0.16523005E-10 0.62476199E+05 0.24622559E+02                   4
C4H2              D11/99C   4H   2    0    0G   300.000  3000.000 1000.        1
 0.91576328E+01 0.55430518E-02-0.13591604E-05 0.18780075E-10 0.23189536E-13    2
 0.52588039E+05-0.23711460E+02 0.10543978E+01 0.41626960E-01-0.65871784E-04    3
 0.53257075E-07-0.16683162E-10 0.54185211E+05 0.14866591E+02                   4
C4H6O25           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
 8.60658242E+00 2.08310051E-02-8.42229481E-06 1.56717640E-09-1.09391202E-13    2
-1.76177415E+04-2.32464750E+01 2.67053463E+00 4.92586420E-03 8.86967406E-05    3
-1.26219194E-07 5.23991321E-11-1.46572472E+04 1.45722395E+01-1.30831522E+04    4
C2H3CHOCH2              C   4H   6O   1    0G   300.000  5000.000 1431.000     1
 1.26762790E+01 1.40819509E-02-4.63473868E-06 7.01090838E-10-3.99438277E-14    2
-4.08065264E+03-4.22515995E+01-3.59388437E+00 5.79063450E-02-4.97163294E-05    3
 2.15818682E-08-3.69199072E-12 8.58852628E+02 4.28475443E+01                   4
C4H4O             T03/97C   4H   4O   1    0G   200.000  6000.0    1000.0      1
 9.38935003E+00 1.40291241E-02-5.07755110E-06 8.24137332E-10-4.95319963E-14    2
-8.68241814E+03-2.79162920E+01 8.47469463E-01 1.31773796E-02 5.99735901E-05    3
-9.71562904E-08 4.22733796E-11-5.36785445E+03 2.14945172E+01-4.17166616E+03    4
C4H6O23           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
 8.60658242E+00 2.08310051E-02-8.42229481E-06 1.56717640E-09-1.09391202E-13    2
-1.32392815E+04-2.32464750E+01 2.67053463E+00 4.92586420E-03 8.86967406E-05    3
-1.26219194E-07 5.23991321E-11-1.02787872E+04 1.45722395E+01-1.30831522E+04    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000     1
 1.39299886E+01 1.13228814E-02-3.87393567E-06 6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01 4.51553480E-01 4.37530418E-02-3.37273602E-05    3
 1.31111496E-08-2.04732021E-12 2.14943141E+03 2.40835867E+01                   4
H2C4O             120189H   2C   4O   1     G  0300.00   4000.00  1000.00      1
 0.01026888E+03 0.04896164E-01-0.04885081E-05-0.02708566E-08 0.05107013E-12    2
 0.02346903E+06-0.02815985E+03 0.04810971E+02 0.01313999E+00 0.09865073E-05    3
-0.06120720E-07 0.01640003E-10 0.02545803E+06 0.02113424E+02                   4
NC3H7CHO   8/12/15      C   4H   8O   1    0G   300.000  5000.000 1679.000     1
 1.19789345E+01 2.04894148E-02-7.24831619E-06 1.15561709E-09-6.84119824E-14    2
-3.09272130E+04-3.63929716E+01 1.24208539E+00 4.21277518E-02-2.13832135E-05    3
 4.22614614E-09-1.03710908E-13-2.71049353E+04 2.21567167E+01                   4
NC3H7CO                 C   4H   7O   1    0G   300.000  5000.000 1496.000     1
 1.34870098E+01 1.58626861E-02-5.41698905E-06 8.40508889E-10-4.87570090E-14    2
-1.30725285E+04-4.38634081E+01 2.63537828E+00 3.40368642E-02-1.24118988E-05    3
-1.17886666E-09 1.16488136E-12-8.65919992E+03 1.68407569E+01                   4
C3H6CHO-1               C   4H   7O   1    0G   300.000  5000.000 1538.000     1
 1.33449137E+01 1.59347421E-02-5.43143577E-06 8.41706117E-10-4.87847084E-14    2
-6.91281947E+03-4.19662475E+01 2.21483383E+00 3.54113290E-02-1.44082892E-05    3
 5.27605922E-11 8.95003230E-13-2.46482792E+03 2.00076022E+01                   4
C3H6CHO-2               C   4H   7O   1    0G   300.000  5000.000 1439.000     1
 1.27128605E+01 1.68632757E-02-5.83779932E-06 9.14059755E-10-5.33575736E-14    2
-8.50165835E+03-3.84620358E+01 4.01372834E+00 2.33173718E-02 5.72463585E-06    3
-1.27182841E-08 3.69912722E-12-4.16766399E+03 1.30545921E+01                   4
C3H6CHO-3               C   4H   7O   1    0G   300.000  5000.000 1678.000     1
 1.21729663E+01 1.80056550E-02-6.43783092E-06 1.03362049E-09-6.14850407E-14    2
-1.08642352E+04-3.80322250E+01 5.29001237E-01 4.30707499E-02-2.49474118E-05    3
 6.40934608E-09-5.27769846E-13-6.87667117E+03 2.48856420E+01                   4
SC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1396.000     1
 1.33892118E+01 1.39115420E-02-4.75820958E-06 7.38736618E-10-4.28606559E-14    2
-1.97917448E+04-4.60146004E+01 1.09372823E+00 4.43315368E-02-3.41918451E-05    3
 1.39369607E-08-2.33791460E-12-1.56745978E+04 1.94458467E+01                   4
SC3H5CO                 C   4H   5O   1    0G   300.000  5000.000 1396.000     1
 1.29925654E+01 1.22140721E-02-4.19305277E-06 6.52697685E-10-3.79407376E-14    2
-2.74782380E+03-4.51092470E+01 7.76401404E-01 4.26828436E-02-3.37881191E-05    3
 1.39128174E-08-2.33331638E-12 1.29903132E+03 1.98102013E+01                   4
C2H5COCH3  8/12/15      C   4H   8O   1    0G   300.000  5000.000 1454.000     1
 1.28183044E+01 1.79874386E-02-5.94194784E-06 9.01636365E-10-5.14993729E-14    2
-3.51711964E+04-4.11609193E+01 2.57048052E+00 3.51446793E-02-1.23849584E-05    3
-1.21280927E-09 1.16163555E-12-3.10194049E+04 1.61395232E+01                   4
C2H5COCH2               C   4H   7O   1    0G   300.000  5000.000 1396.000     1
 1.35979480E+01 1.57187785E-02-5.35200820E-06 8.28428039E-10-4.79645862E-14    2
-1.30111973E+04-4.46215708E+01 1.96643032E+00 4.10271409E-02-2.56193885E-05    3
 7.86244495E-09-9.26825962E-13-8.80149212E+03 1.84803948E+01                   4
CH2CH2COCH3             C   4H   7O   1    0G   300.000  5000.000 1392.000     1
 1.17915603E+01 1.70296457E-02-5.75444256E-06 8.86035114E-10-5.11070778E-14    2
-9.70683178E+03-3.25532787E+01 2.36191763E+00 3.50400641E-02-1.70487065E-05    3
 3.09070210E-09 2.80364847E-14-6.02754073E+03 1.95184512E+01                   4
CH3CHCOCH3              C   4H   7O   1    0G   300.000  5000.000 1438.000     1
 1.19651378E+01 1.63142163E-02-5.39879520E-06 8.20454677E-10-4.69197541E-14    2
-1.51990676E+04-3.30142593E+01 3.31082456E+00 2.83712402E-02-5.64603859E-06    3
-4.62626296E-09 1.82954207E-12-1.14602301E+04 1.62217415E+01                   4
C2H3COCH3               C   4H   6O   1    0G   300.000  5000.000 1390.000     1
 1.19989844E+01 1.52616304E-02-5.26018882E-06 8.20774274E-10-4.77834528E-14    2
-2.12170620E+04-3.71383523E+01 6.55910700E-01 4.19405303E-02-3.00269693E-05    3
 1.16578089E-08-1.92100897E-12-1.72216627E+04 2.38412293E+01                   4
CH3CHOOCOCH3            C   4H   7O   3    0G   300.000  5000.000 1411.000     1
 1.68056216E+01 1.70791389E-02-5.69439450E-06 8.68878944E-10-4.98008338E-14    2
-3.06718613E+04-5.51178960E+01 4.30171569E+00 4.62273591E-02-3.12564494E-05    3
 1.08627824E-08-1.51478379E-12-2.63732146E+04 1.19724375E+01                   4
CH2CHOOHCOCH3           C   4H   7O   3    0G   300.000  5000.000 1413.000     1
 1.78031394E+01 1.60286227E-02-5.38152372E-06 8.25242310E-10-4.74718968E-14    2
-2.30767899E+04-5.87370258E+01 4.45962223E+00 4.67200276E-02-3.15878907E-05    3
 1.06245787E-08-1.38857032E-12-1.84720686E+04 1.29655977E+01                   4
C2H5CHCO                C   4H   6O   1    0G   300.000  5000.000 1550.000     1
-2.04040652E+02 2.93466880E-01-1.15884523E-04 1.95253673E-08-1.19030791E-12    2
 8.27380036E+04 1.21233386E+03-2.28307043E+01 1.70978191E-01-3.53394379E-04    3
 2.78221616E-07-6.77325074E-11-1.04125457E+04 1.31232921E+02                   4
IC4H6Q2-II 9/ 8/14      C   4H   8O   4    0G   300.000  5000.000 1386.000     1
 2.50360805E+01 1.60230197E-02-5.70704966E-06 9.10412038E-10-5.38294659E-14    2
-2.84196401E+04-9.67186452E+01 2.16408482E-01 8.25572149E-02-7.64540445E-05    3
 3.58211787E-08-6.67718658E-12-2.05694845E+04 3.36943223E+01                   4
C5H10-1                 C   5H  10    0    0G   300.000  5000.000 1390.000     1
 1.43624894E+01 2.26076154E-02-7.70500843E-06 1.19329968E-09-6.91126022E-14    2
-9.99915627E+03-5.12512094E+01-1.65023816E-01 5.30727359E-02-3.10861587E-05    3
 8.92413402E-09-9.81619602E-13-4.57363143E+03 2.80570113E+01                   4
C5H81-3    9/ 8/14      C   5H   8    0    0G   300.000  5000.000 1385.000     1
 1.29945372E+01 1.92678312E-02-6.58966712E-06 1.02295969E-09-5.93441369E-14    2
 4.59040047E+03-4.35689825E+01 1.54882436E+00 4.15042709E-02-2.14359890E-05    3
 4.71145517E-09-2.42142508E-13 9.05636062E+03 1.95665910E+01                   4
C5H9O1-3   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1379.000     1
 1.78860333E+01 2.04837367E-02-7.16613461E-06 1.12948597E-09-6.62221468E-14    2
-4.33139568E+03-6.72851315E+01 2.49666166E+00 5.20326105E-02-3.09828268E-05    3
 9.02567482E-09-1.04311127E-12 1.54758549E+03 1.70868328E+01                   4
BC5H10     9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1389.000     1
 1.40426423E+01 2.27915348E-02-7.74902598E-06 1.19814522E-09-6.93127003E-14    2
-1.32160483E+04-5.14469569E+01 6.04882839E-01 4.96635256E-02-2.66571142E-05    3
 6.47312078E-09-4.84017883E-13-8.06312207E+03 2.23818263E+01                   4
CC5H9-A                 C   5H   9    0    0G   300.000  5000.000 1393.000     1
 1.38635892E+01 2.06362872E-02-7.05717373E-06 1.09539676E-09-6.35381849E-14    2
 1.36104251E+04-4.72507189E+01-6.78909715E-01 5.37496002E-02-3.61116825E-05    3
 1.28563411E-08-1.92155723E-12 1.87974429E+04 3.12403382E+01                   4
CC5H9-B    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1392.000     1
 1.35249511E+01 2.14363755E-02-7.35304116E-06 1.14368637E-09-6.64363518E-14    2
 5.41381916E+03-5.00302394E+01-6.91501860E-01 5.09804846E-02-2.96448293E-05    3
 8.28273022E-09-8.57575066E-13 1.07478467E+04 2.76711552E+01                   4
AC5H9O-C                C   5H   9O   1    0G   300.000  5000.000 1382.000     1
 1.76789601E+01 2.05915073E-02-7.18764438E-06 1.13116483E-09-6.62505034E-14    2
-6.25146818E+03-6.62131721E+01 2.04951318E+00 5.36584877E-02-3.35086710E-05    3
 1.06174235E-08-1.39224338E-12-3.85112518E+02 1.91077262E+01                   4
CC5H9O-B   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1377.000     1
 1.86974377E+01 1.84542537E-02-6.18682537E-06 9.48850967E-10-5.46203980E-14    2
-7.15897769E+03-7.26540429E+01 2.75614808E+00 5.20514036E-02-3.10966938E-05    3
 8.25895065E-09-6.59917121E-13-1.35162741E+03 1.40990119E+01                   4
AC5H10                  C   5H  10    0    0G   300.000  5000.000 1392.000     1
 1.41931279E+01 2.26551019E-02-7.70008627E-06 1.19031326E-09-6.88489604E-14    2
-1.19491010E+04-5.10688681E+01-5.39429136E-01 5.44489715E-02-3.32707895E-05    3
 1.03047694E-08-1.28363329E-12-6.53967251E+03 2.90349986E+01                   4
AC5H9-A2                C   5H   9    0    0G   300.000  5000.000 1385.000     1
 1.50019889E+01 1.95965428E-02-6.60205927E-06 1.01535593E-09-5.85454957E-14    2
 5.90081014E+03-5.54528992E+01-9.54047710E-01 5.50153471E-02-3.58307910E-05    3
 1.16444141E-08-1.49086833E-12 1.15959514E+04 3.08476806E+01                   4
AC5H9-C                 C   5H   9    0    0G   300.000  5000.000 1392.000     1
 1.37918110E+01 2.09644966E-02-7.13793293E-06 1.10480881E-09-6.39628018E-14    2
 5.09555600E+03-5.01391436E+01-8.41372657E-01 5.27157283E-02-3.27334707E-05    3
 1.01974035E-08-1.26084730E-12 1.04321036E+04 2.93316754E+01                   4
AC5H9-D                 C   5H   9    0    0G   300.000  5000.000 1393.000     1
 1.35607521E+01 2.07514878E-02-7.06608626E-06 1.09362345E-09-6.33083050E-14    2
 1.31896844E+04-4.48718988E+01-1.67398152E-01 5.09876974E-02-3.22615638E-05    3
 1.05911843E-08-1.43705463E-12 1.81792947E+04 2.95710715E+01                   4
B2E2M1OJ                C   5H   9O   1    0G   300.000  5000.000 2003.000     1
 1.35666458E+01 2.56547934E-02-9.37226256E-06 1.52518398E-09-9.15378763E-14    2
-3.58767067E+03-4.27272791E+01 5.64762692E+00 3.43609862E-02-5.60649548E-06    3
-5.19111402E-09 1.73155461E-12-6.65737793E+00 3.13825267E+00                   4
B13DE2M                 C   5H   8    0    0G   300.000  5000.000 1397.000     1
 1.40757545E+01 1.82375566E-02-6.20747687E-06 9.60350919E-10-5.55741525E-14    2
 2.40033881E+03-5.12988284E+01-4.72170009E-01 5.59413257E-02-4.50458826E-05    3
 1.96181377E-08-3.52009647E-12 7.14960489E+03 2.56276807E+01                   4
B13DE2MJ                C   5H   7    0    0G   300.000  5000.000 1393.000     1
 1.48413344E+01 1.52425753E-02-5.13559858E-06 7.89787260E-10-4.55353492E-14    2
 2.02661570E+04-5.54474955E+01-8.98037227E-01 5.65174321E-02-4.76107829E-05    3
 2.09672106E-08-3.73076319E-12 2.52881763E+04 2.74966602E+01                   4
B12DE3M   11/12/12 THERMC   5H   8    0    0G   300.000  5000.000 1388.000     1
 1.37093177E+01 1.85726726E-02-6.33115904E-06 9.80719059E-10-5.68099894E-14    2
 8.59518752E+03-4.88749621E+01 1.27860173E+00 4.54917474E-02-2.82334169E-05    3
 8.98449372E-09-1.17220042E-12 1.31637341E+04 1.87039373E+01                   4
B2E3M1OJ                C   5H   9O   1    0G   300.000  5000.000 2003.000     1
 1.35666458E+01 2.56547934E-02-9.37226256E-06 1.52518398E-09-9.15378763E-14    2
-3.58767067E+03-4.27272791E+01 5.64762692E+00 3.43609862E-02-5.60649548E-06    3
-5.19111402E-09 1.73155461E-12-6.65737793E+00 3.13825267E+00                   4
TC4H8CHO   9/ 7/95 THERMC   5H   9O   1    0G   300.000  5000.000 1397.00      1
 1.79663933E+01 1.94207117E-02-6.67409451E-06 1.03969221E-09-6.04702651E-14    2
-1.33368585E+04-6.79819424E+01-9.58078294E-01 6.42003258E-02-4.70776827E-05    3
 1.75737698E-08-2.64896151E-12-6.86582501E+03 3.33781112E+01                   4
O2C4H8CHO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1395.00      1
 2.12629904E+01 2.14072282E-02-7.38342949E-06 1.15281523E-09-6.71508438E-14    2
-3.16854524E+04-7.99828703E+01 1.91847699E+00 6.67245869E-02-4.80871046E-05    3
 1.78588690E-08-2.71163880E-12-2.49837984E+04 2.38577867E+01                   4
O2HC4H8CO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1394.00      1
 2.38219630E+01 1.91411448E-02-6.67919154E-06 1.05127303E-09-6.15876805E-14    2
-3.23093973E+04-9.42580755E+01 1.82607262E+00 6.93466111E-02-4.93125140E-05    3
 1.69848340E-08-2.26117657E-12-2.46578311E+04 2.41167544E+01                   4
C6H101-5   4/12/13 THERMC   6H  10    0    0G   300.000  5000.000 1413.000     1
 1.60456030E+01 2.34774145E-02-7.85797929E-06 1.20200542E-09-6.90100029E-14    2
 2.11899382E+03-5.88452460E+01-1.01375402E+00 6.38242808E-02-4.40653860E-05    3
 1.58295163E-08-2.30830701E-12 7.94033696E+03 3.25056094E+01                   4
C6H9-A    12/ 5/12 THERMC   6H   9    0    0G   300.000  5000.000 1400.000     1
 1.70842767E+01 2.08842788E-02-7.14529004E-06 1.10943563E-09-6.43676989E-14    2
 2.01040204E+04-6.39326012E+01-2.66715213E+00 7.26196475E-02-6.05323920E-05    3
 2.66000571E-08-4.74613408E-12 2.64415017E+04 4.02220332E+01                   4
H15DE25DM               C   8H  14    0    0G   300.000  5000.000 1395.000     1
 2.25355644E+01 3.23955734E-02-1.10270814E-05 1.70640907E-09-9.87758061E-14    2
-1.04808866E+04-9.19784905E+01-1.71853441E+00 8.82613783E-02-6.03140500E-05    3
 2.15862289E-08-3.19690882E-12-1.95255748E+03 3.86048681E+01                   4
H15DE25DM-S             C   8H  13    0    0G   300.000  5000.000 1395.000     1
 2.21422958E+01 3.06966055E-02-1.04617380E-05 1.62037747E-09-9.38578511E-14    2
 6.56045671E+03-9.04059585E+01-2.04235551E+00 8.66261688E-02-5.99110976E-05    3
 2.15551630E-08-3.18976697E-12 1.50224279E+04 3.96917763E+01                   4
H15DE25DM-A             C   8H  13    0    0G   300.000  5000.000 1391.000     1
 2.33282646E+01 2.93694154E-02-9.94258906E-06 1.53368063E-09-8.86030202E-14    2
 7.37319036E+03-9.55902415E+01-2.21863377E+00 8.91652629E-02-6.33360636E-05    3
 2.32007379E-08-3.46329567E-12 1.61971179E+04 4.15116620E+01                   4
H15DE25DM-AO            C   8H  13O   1    0G   300.000  5000.000 1378.000     1
 2.50985951E+01 3.15085628E-02-1.10076915E-05 1.73332426E-09-1.01557468E-13    2
-2.49465338E+03-1.01097942E+02 3.03691957E+00 7.50640438E-02-4.17779534E-05    3
 1.07915725E-08-9.97734397E-13 6.11649780E+03 2.04746031E+01                   4
H15DE25DM-SO            C   8H  13O   1    0G   300.000  5000.000 1388.000     1
 2.60152179E+01 3.04295766E-02-1.05676513E-05 1.65746547E-09-9.68470091E-14    2
-4.79568520E+03-1.06442472E+02 9.30464015E-01 8.71669873E-02-5.99582593E-05    3
 2.15026041E-08-3.21687573E-12 4.19310073E+03 2.90924508E+01                   4
H15DE2M-T               C   7H  11    0    0G   300.000  5000.000 1389.000     1
 1.90144729E+01 2.61932198E-02-9.01183878E-06 1.40455988E-09-8.17075251E-14    2
 2.35551101E+04-7.15568628E+01 3.88856066E-01 6.70215700E-02-4.29671268E-05    3
 1.42489875E-08-1.96105571E-12 3.03627273E+04 2.95444186E+01                   4
IC4H7CHO                C   5H   8O   1    0G   300.000  5000.000 1391.000     1
 1.59171638E+01 1.93357284E-02-6.70857943E-06 1.05155191E-09-6.14175906E-14    2
-2.16140735E+04-5.67616631E+01-1.20982776E+00 5.92603375E-02-4.26960089E-05    3
 1.60356164E-08-2.49347521E-12-1.56205327E+04 3.53137305E+01                   4
L-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
 0.12715182E+02 0.13839662E-01-0.43765440E-05 0.31541636E-09 0.46619026E-13    2
 0.57031148E+05-0.39464600E+02 0.29590225E+00 0.58053318E-01-0.67766756E-04    3
 0.43376762E-07-0.11418864E-10 0.60001371E+05 0.22318970E+02                   4
C-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
 0.13849209E+02 0.78807920E-02 0.18243836E-05-0.21169166E-08 0.37459977E-12    2
 0.47446340E+05-0.50404953E+02-0.30991268E+01 0.54030564E-01-0.40839004E-04    3
 0.10738837E-07 0.98078490E-12 0.52205711E+05 0.37415207E+02                   4
C6H3              H6W/94C   6H   3    0    0G   300.000  3000.00  1000.00      1
 0.58188343E+01 0.27933408E-01-0.17825427E-04 0.53702536E-08-0.61707627E-12    2
 0.85188250E+05-0.92147827E+00 0.11790619E+01 0.55547360E-01-0.73076168E-04    3
 0.52076736E-07-0.15046964E-10 0.85647312E+05 0.19179199E+02                   4
C6H2              P 1/93C   6H   2    0    0G   300.000  3000.00  1000.00      1
 0.13226281E+02 0.73904302E-02-0.22715381E-05 0.25875217E-09-0.55356741E-14    2
 0.80565258E+05-0.41201176E+02-0.15932624E+01 0.80530145E-01-0.14800649E-03    3
 0.13300031E-06-0.45332313E-10 0.83273227E+05 0.27980873E+02                   4
C6H6              G 6/01C   6H   6    0    0G   200.000  6000.000 1000.000     1
 1.10809576E+01 2.07176746E-02-7.52145991E-06 1.22320984E-09-7.36091279E-14    2
 4.30641035E+03-4.00413310E+01 5.04818632E-01 1.85020642E-02 7.38345881E-05    3
-1.18135741E-07 5.07210429E-11 8.55247913E+03 2.16412893E+01 9.96811598E+03    4
FULVENE                0C   6H   6    0    0G   200.000  5000.000 1000.00      1
 0.11103525E+02 0.20600685E-01-0.75302224E-05 0.12388695E-08-0.75415976E-13    2
 0.20361843E+05-0.36665197E+02-0.71813191E+00 0.37934312E-01 0.11398837E-04    3
-0.41333503E-07 0.18055927E-10 0.24223825E+05 0.27855714E+02                   4
C6H5              T04/02C   6H   5    0    0G   200.000  6000.000 1000.        1
 1.08444762E+01 1.73212473E-02-6.29233249E-06 1.02369961E-09-6.16216828E-14    2
 3.55598475E+04-3.53735134E+01 2.10306633E-01 2.04745507E-02 5.89743006E-05    3
-1.01534255E-07 4.47105660E-11 3.95468722E+04 2.52910455E+01 4.08610970E+04    4
C6H5OO     3/26/ 9 THERMC   6H   5O   2    0G   300.000  5000.000 1403.000     1
 1.67078262E+01 1.62326229E-02-5.47969630E-06 8.43510060E-10-4.86562431E-14    2
 8.14242915E+03-6.08346973E+01-2.99164672E+00 7.03857150E-02-6.34400574E-05    3
 2.91548920E-08-5.30706938E-12 1.41320240E+04 4.20142955E+01                   4
C6H5OOH    3/26/ 9 THERMC   6H   6O   2    0G   300.000  5000.000 1404.000     1
 1.92317474E+01 1.63154699E-02-5.53448904E-06 8.55059974E-10-4.94583790E-14    2
-1.01971012E+04-7.61674471E+01-4.03105975E+00 7.96101888E-02-7.21655013E-05    3
 3.27610696E-08-5.85584239E-12-3.10973017E+03 4.54324978E+01                   4
C6H5OH            L 4/84C   6H   6O   1    0G   300.000  5000.000 1000.        1
 0.14912073E+02 0.18378135E-01-0.61983128E-05 0.91983221E-09-0.49209565E-13    2
-0.18375199E+05-0.55924103E+02-0.16956539E+01 0.52271299E-01-0.72024050E-05    3
-0.35859603E-07 0.20449073E-10-0.13284121E+05 0.32542160E+02-0.11594207E+05    4
C6H5O             T05/02C   6H   5O   1    0G   200.000  6000.000 1000.        1
 1.37221720E+01 1.74688771E-02-6.35504520E-06 1.03492308E-09-6.23410504E-14    2
 2.87274751E+02-4.88181680E+01-4.66204455E-01 4.13443975E-02 1.32412991E-05    3
-5.72872769E-08 2.89763707E-11 4.77858391E+03 2.76990274E+01 6.49467016E+03    4
C6H4OH     4/ 9/ 9 THERMC   6H   5O   1    0G   300.000  5000.000 1402.000     1
 1.73187560E+01 1.36366984E-02-4.68316332E-06 7.29071204E-10-4.23805358E-14    2
 1.14990276E+04-6.89986593E+01-5.99875435E+00 8.59063379E-02-9.12525636E-05    3
 4.72275890E-08-9.35576749E-12 1.78621926E+04 4.99931427E+01                   4
OC6H4OH    4/ 9/ 9 THERMC   6H   5O   2    0G   300.000  5000.000 1403.000     1
 2.22718210E+01 1.21038561E-02-4.18429526E-06 6.54475399E-10-3.81746504E-14    2
-2.34827539E+04-9.61035467E+01-8.02205657E+00 1.09403210E-01-1.23489276E-04    3
 6.56286805E-08-1.31527870E-11-1.55949156E+04 5.72175202E+01                   4
O-C6H4O2          AK0405C   6H   4O   2    0G   270.000  3000.000 1370.00      1
 1.23614349E+01 2.40491397E-02-1.16529057E-05 2.71332785E-09-2.47593219E-13    2
-1.67079717E+04-4.00310857E+01-2.36179712E+00 6.86058343E-02-6.39129516E-05    3
 3.06903009E-08-5.97357785E-12-1.26704431E+04 3.53724482E+01                   4
P-C6H4O2          AK0405C   6H   4O   2    0G   270.000  3000.000 1370.00      1
 1.23423732E+01 2.40612690E-02-1.16565184E-05 2.71393504E-09-2.47643065E-13    2
-2.06185312E+04-4.08244024E+01-2.43170113E+00 6.87937608E-02-6.41382837E-05    3
 3.08126855E-08-5.99832072E-12-1.65696994E+04 3.48309430E+01                   4
O-OC6H5OJ  WKM          C   6O   2H   5    0G   300.000  5000.000 1400.000     1
 1.84625733E+01 1.57607263E-02-5.44671499E-06 8.51765760E-10-4.96759541E-14    2
-1.72770226E+02-7.28742484E+01-2.65459198E+00 7.17179095E-02-6.31552372E-05    3
 2.81132946E-08-4.97463333E-12 6.45283150E+03 3.81123139E+01                   4
P-OC6H5OJ  WKM          C   6O   2H   5    0G   300.000  5000.000 1400.000     1
 1.82799770E+01 1.59280974E-02-5.50765220E-06 8.61649836E-10-5.02677539E-14    2
-6.25907994E+01-7.25809444E+01-3.29683290E+00 7.27365977E-02-6.36158220E-05    3
 2.80683553E-08-4.92279426E-12 6.73402222E+03 4.09349895E+01                   4
P-C6H3O2          AK0505C   6H   3O   2    0G   270.000  3000.000 1290.00      1
 1.22963699E+01 2.15055142E-02-1.07516136E-05 2.57528163E-09-2.41023652E-13    2
 1.15428998E+04-3.72584002E+01-1.57852347E+00 6.55376473E-02-6.50308721E-05    3
 3.32026554E-08-6.86665555E-12 1.51750093E+04 3.31518638E+01                   4
C5H6              T 1/90C   5H   6    0    0G   200.000  6000.000 1000.        1
 0.99757848E+01 0.18905543E-01-0.68411461E-05 0.11099340E-08-0.66680236E-13    2
 0.11081693E+05-0.32209454E+02 0.86108957E+00 0.14804031E-01 0.72108895E-04    3
-0.11338055E-06 0.48689972E-10 0.14801755E+05 0.21353453E+02 0.16152485E+05    4
C5H5             TAK0505C   5H   5    0    0G   298.150  3500.000  969.35      1
 1.33675715E+00 3.24793912E-02-1.67587774E-05 4.03514137E-09-3.70739036E-13    2
 3.00730524E+04 1.60315806E+01-3.97555452E+00 7.41370991E-02-1.11803345E-04    3
 9.04628776E-08-2.80999747E-11 3.01769405E+04 3.67153636E+01                   4
C5H6-L     2/ 5/ 9 THERMC   5H   6    0    0G   300.000  5000.000 1372.000     1
 1.29600892E+01 1.48953758E-02-5.23622902E-06 8.27916389E-10-4.86464523E-14    2
 2.38180800E+04-4.25312093E+01 3.58448213E+00 3.24459626E-02-1.70150991E-05    3
 4.22715914E-09-4.18452556E-13 2.76514681E+04 9.60644208E+00                   4
C#CCVCCJ           GLAR C   5H   5    0    0G   300.000  5000.000 1396.000     1
 1.41230912E+01 1.14233190E-02-3.95851276E-06 6.20128961E-10-3.62097887E-14    2
 4.25158384E+04-5.02942871E+01-6.16143558E-01 5.06466579E-02-4.48561743E-05    3
 2.02459419E-08-3.64542145E-12 4.71532377E+04 2.71623299E+01                   4
C5H7       1/22/ 9 WKM  C   5H   7    0    0G   300.000  5000.000 1377.000     1
 1.36630213E+01 1.68061358E-02-5.98746539E-06 9.55341072E-10-5.64951981E-14    2
 1.27238941E+04-5.46331286E+01-6.75118368E+00 6.06461693E-02-4.01260152E-05    3
 1.22051562E-08-1.33459844E-12 2.01365277E+04 5.62694938E+01                   4
CVCCJCVC   3/1/95  Z&B  C   5H   7    0    0G   300.000  5000.000 1388.000     1
 1.40879309E+01 1.62398907E-02-5.64768950E-06 8.86857524E-10-5.18698993E-14    2
 1.76798698E+04-5.13735038E+01-2.94595603E+00 5.68783623E-02-4.31336497E-05    3
 1.68169537E-08-2.67926433E-12 2.35156925E+04 3.98188778E+01                   4
CVCCVCCJ           Z&B  C   5H   7    0    0G   300.000  5000.000 1386.000     1
 1.47302883E+01 1.59030900E-02-5.57729508E-06 8.80604825E-10-5.16963733E-14    2
 1.74050791E+04-5.42670706E+01-1.60087476E+00 5.38764703E-02-3.96302225E-05    3
 1.49599474E-08-2.31995284E-12 2.31199746E+04 3.35492960E+01                   4
CVCCJCVCOH 10/6/95 Z&B  C   5H   7O   1    0G   300.000  5000.000 1397.000     1
 1.67465815E+01 1.58357240E-02-5.44954706E-06 8.49881387E-10-4.94743246E-14    2
-4.30972870E+03-6.19378748E+01-2.91175436E+00 6.69362484E-02-5.71603047E-05    3
 2.48753749E-08-4.33243894E-12 1.96441523E+03 4.17454344E+01                   4
HOCVCCVO   1/26/ 9 WKM  C   3H   4O   2    0G   300.000  5000.000 1413.000     1
 1.66505478E+01 6.11745137E-03-2.09080785E-06 3.24985683E-10-1.88875073E-14    2
-3.82179939E+04-6.36794754E+01-2.01837189E+00 6.26539783E-02-6.73359280E-05    3
 3.39430425E-08-6.48917648E-12-3.31367523E+04 3.18162860E+01                   4
CVCCVCCOH  1/23/ 9 WKM  C   5H   8O   1    0G   300.000  5000.000 1396.000     1
 1.63079670E+01 1.79957763E-02-6.03115896E-06 9.23992259E-10-5.31254053E-14    2
-1.58204603E+04-5.84137244E+01-5.31488384E-01 6.06983915E-02-4.81499862E-05    3
 2.00308244E-08-3.38987282E-12-1.03301302E+04 3.07961436E+01                   4
OC5H7O     1/22/ 9 WKM  C   5H   7O   2    0G   300.000  5000.000 1375.000     1
 1.65416953E+01 1.86677673E-02-6.44836048E-06 1.00787611E-09-5.87521858E-14    2
-2.82017168E+04-5.47258181E+01 4.88394767E+00 4.03401300E-02-1.97774150E-05    3
 3.68903501E-09-3.40202384E-14-2.35295942E+04 9.97070337E+00                   4
OC4H6O     1/23/ 9 WKM  C   4H   6O   2    0G   300.000  5000.000 1382.000     1
 1.41894774E+01 1.53345510E-02-5.24594862E-06 8.14655154E-10-4.72759368E-14    2
-4.10001835E+04-4.43771751E+01 4.21628848E+00 3.57422725E-02-2.04226185E-05    3
 5.63821367E-09-5.88888993E-13-3.72055911E+04 1.02814620E+01                   4
OC4H5O     1/23/ 9 WKM  C   4H   5O   2    0G   300.000  5000.000 1388.000     1
 1.32138775E+01 1.37339051E-02-4.62639517E-06 7.10941370E-10-4.09538499E-14    2
-2.16535271E+04-3.64185255E+01 4.60550978E+00 3.30498712E-02-2.13102363E-05    3
 7.37021089E-09-1.08289438E-12-1.85460831E+04 1.01599453E+01                   4
O2CCHOOJ           Z&B  C   2H   1O   4    0G   300.000  5000.000 1682.000     1
 1.09910849E+01 7.46985861E-03-2.75568271E-06 4.51353051E-10-2.72108652E-14    2
-3.51335323E+04-2.11652231E+01 8.91497688E+00 8.60571847E-03 5.24416766E-07    3
-2.79301331E-09 7.62963051E-13-3.40867754E+04-8.72978273E+00                   4
HOCVCCJVO  1/26/ 9 WKM  C   3H   3O   2    0G   300.000  5000.000 1414.000     1
 1.52720985E+01 5.02586331E-03-1.68408578E-06 2.58390706E-10-1.48849424E-14    2
-1.98506828E+04-5.54641734E+01 6.07270082E-01 4.96011303E-02-5.32300885E-05    3
 2.68392951E-08-5.13094510E-12-1.58814562E+04 1.94817133E+01                   4
C5H5OH     5/ 2/91 THE.MC   5H   6O   1    0G   300.000  5000.000 1398.000     1
 1.53433477E+01 1.50754059E-02-5.13553582E-06 7.95807816E-10-4.61311517E-14    2
-1.19645453E+04-5.85204430E+01-4.26822012E+00 6.62446749E-02-5.68494038E-05    3
 2.46858526E-08-4.26820696E-12-5.75581338E+03 4.47962850E+01                   4
C5H5O      5/16/90 THERMC   5H   5O   1    0G   300.000  5000.000 1392.000     1
 1.48322894E+01 1.40483376E-02-4.92302051E-06 7.77041219E-10-4.56103939E-14    2
 1.45523665E+04-5.73228191E+01-2.83112840E+00 5.67277287E-02-4.44757303E-05    3
 1.74924447E-08-2.76004847E-12 2.04992154E+04 3.69634411E+01                   4
C5H4OH            T 8/99C   5H   5O   1    0G   200.000  6000.000 1000.        1
 1.33741248E+01 1.51996469E-02-5.45685046E-06 8.80944866E-10-5.27493258E-14    2
 2.20358027E+03-4.59569069E+01-1.28398054E+00 4.90298511E-02-1.35844414E-05    3
-2.92983743E-08 1.90820619E-11 6.37364803E+03 3.08073591E+01 8.00114499E+03    4
C5H4O             T 8/99C   5H   4O   1    0G   200.000  6000.000 1000.        1
 1.00806824E+01 1.61143465E-02-5.83314509E-06 9.46759320E-10-5.68972206E-14    2
 1.94364771E+03-2.94521623E+01 2.64576497E-01 3.34873827E-02 1.67738470E-06    3
-2.96207455E-08 1.54431476E-11 5.11159287E+03 2.35409513E+01 6.64245999E+03    4
C5H3O            TAK0905C   5H   3O   1    0G   300.000  3500.000 1500.00      1
 1.19961781E+01 1.34287065E-02-5.90045309E-06 1.22553862E-09-9.86114716E-14    2
 2.89592010E+04-4.07548249E+01-3.03242604E+00 5.43937201E-02-4.95018348E-05    3
 2.25523751E-08-4.10727920E-12 3.35644081E+04 3.78374823E+01                   4
CJVCCVCCVO 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1396.000     1
 1.62360823E+01 1.18297101E-02-4.11454219E-06 6.46026823E-10-3.77767639E-14    2
 1.93499885E+04-5.83498817E+01-5.06628841E-01 6.04671965E-02-5.97396749E-05    3
 2.96804228E-08-5.76240010E-12 2.42765544E+04 2.82994148E+01                   4
CVCCVCCJVO 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1399.000     1
 1.53178248E+01 1.27352911E-02-4.35882964E-06 6.76912763E-10-3.92771371E-14    2
 7.60582726E+03-5.43599625E+01-2.18492198E-01 5.92100223E-02-5.89241174E-05    3
 2.97411920E-08-5.85244770E-12 1.20600764E+04 2.55968530E+01                   4
CJVCCVO    4/ 8/94 THERMC   3H   3O   1    0G   300.000  5000.000 1402.000     1
 1.07482537E+01 6.19822688E-03-2.06130981E-06 3.14418872E-10-1.80309517E-14    2
 1.51410162E+04-3.01266033E+01 1.46654466E+00 3.23390476E-02-3.05588208E-05    3
 1.44081861E-08-2.65600505E-12 1.78850058E+04 1.80850321E+01                   4
END
